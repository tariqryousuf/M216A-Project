module pix_mem(
	input clk,
	input enable,
	input [9:0]  Pix_0, Pix_1, Pix_2, Pix_3, Pix_4, Pix_5, Pix_6, Pix_7, Pix_8, Pix_9, Pix_10, Pix_11, Pix_12, Pix_13, Pix_14, Pix_15, Pix_16, Pix_17, Pix_18, Pix_19, Pix_20, Pix_21, Pix_22, Pix_23, Pix_24, Pix_25, Pix_26, Pix_27, Pix_28, Pix_29, Pix_30, Pix_31, Pix_32, Pix_33, Pix_34, Pix_35, Pix_36, Pix_37, Pix_38, Pix_39, Pix_40, Pix_41, Pix_42, Pix_43, Pix_44, Pix_45, Pix_46, Pix_47, Pix_48, Pix_49, Pix_50, Pix_51, Pix_52, Pix_53, Pix_54, Pix_55, Pix_56, Pix_57, Pix_58, Pix_59, Pix_60, Pix_61, Pix_62, Pix_63, Pix_64, Pix_65, Pix_66, Pix_67, Pix_68, Pix_69, Pix_70, Pix_71, Pix_72, Pix_73, Pix_74, Pix_75, Pix_76, Pix_77, Pix_78, Pix_79, Pix_80, Pix_81, Pix_82, Pix_83, Pix_84, Pix_85, Pix_86, Pix_87, Pix_88, Pix_89, Pix_90, Pix_91, Pix_92, Pix_93, Pix_94, Pix_95, Pix_96, Pix_97, Pix_98, Pix_99, Pix_100, Pix_101, Pix_102, Pix_103, Pix_104, Pix_105, Pix_106, Pix_107, Pix_108, Pix_109, Pix_110, Pix_111, Pix_112, Pix_113, Pix_114, Pix_115, Pix_116, Pix_117, Pix_118, Pix_119, Pix_120, Pix_121, Pix_122, Pix_123, Pix_124, Pix_125, Pix_126, Pix_127, Pix_128, Pix_129, Pix_130, Pix_131, Pix_132, Pix_133, Pix_134, Pix_135, Pix_136, Pix_137, Pix_138, Pix_139, Pix_140, Pix_141, Pix_142, Pix_143, Pix_144, Pix_145, Pix_146, Pix_147, Pix_148, Pix_149, Pix_150, Pix_151, Pix_152, Pix_153, Pix_154, Pix_155, Pix_156, Pix_157, Pix_158, Pix_159, Pix_160, Pix_161, Pix_162, Pix_163, Pix_164, Pix_165, Pix_166, Pix_167, Pix_168, Pix_169, Pix_170, Pix_171, Pix_172, Pix_173, Pix_174, Pix_175, Pix_176, Pix_177, Pix_178, Pix_179, Pix_180, Pix_181, Pix_182, Pix_183, Pix_184, Pix_185, Pix_186, Pix_187, Pix_188, Pix_189, Pix_190, Pix_191, Pix_192, Pix_193, Pix_194, Pix_195, Pix_196, Pix_197, Pix_198, Pix_199, Pix_200, Pix_201, Pix_202, Pix_203, Pix_204, Pix_205, Pix_206, Pix_207, Pix_208, Pix_209, Pix_210, Pix_211, Pix_212, Pix_213, Pix_214, Pix_215, Pix_216, Pix_217, Pix_218, Pix_219, Pix_220, Pix_221, Pix_222, Pix_223, Pix_224, Pix_225, Pix_226, Pix_227, Pix_228, Pix_229, Pix_230, Pix_231, Pix_232, Pix_233, Pix_234, Pix_235, Pix_236, Pix_237, Pix_238, Pix_239, Pix_240, Pix_241, Pix_242, Pix_243, Pix_244, Pix_245, Pix_246, Pix_247, Pix_248, Pix_249, Pix_250, Pix_251, Pix_252, Pix_253, Pix_254, Pix_255, Pix_256, Pix_257, Pix_258, Pix_259, Pix_260, Pix_261, Pix_262, Pix_263, Pix_264, Pix_265, Pix_266, Pix_267, Pix_268, Pix_269, Pix_270, Pix_271, Pix_272, Pix_273, Pix_274, Pix_275, Pix_276, Pix_277, Pix_278, Pix_279, Pix_280, Pix_281, Pix_282, Pix_283, Pix_284, Pix_285, Pix_286, Pix_287, Pix_288, Pix_289, Pix_290, Pix_291, Pix_292, Pix_293, Pix_294, Pix_295, Pix_296, Pix_297, Pix_298, Pix_299, Pix_300, Pix_301, Pix_302, Pix_303, Pix_304, Pix_305, Pix_306, Pix_307, Pix_308, Pix_309, Pix_310, Pix_311, Pix_312, Pix_313, Pix_314, Pix_315, Pix_316, Pix_317, Pix_318, Pix_319, Pix_320, Pix_321, Pix_322, Pix_323, Pix_324, Pix_325, Pix_326, Pix_327, Pix_328, Pix_329, Pix_330, Pix_331, Pix_332, Pix_333, Pix_334, Pix_335, Pix_336, Pix_337, Pix_338, Pix_339, Pix_340, Pix_341, Pix_342, Pix_343, Pix_344, Pix_345, Pix_346, Pix_347, Pix_348, Pix_349, Pix_350, Pix_351, Pix_352, Pix_353, Pix_354, Pix_355, Pix_356, Pix_357, Pix_358, Pix_359, Pix_360, Pix_361, Pix_362, Pix_363, Pix_364, Pix_365, Pix_366, Pix_367, Pix_368, Pix_369, Pix_370, Pix_371, Pix_372, Pix_373, Pix_374, Pix_375, Pix_376, Pix_377, Pix_378, Pix_379, Pix_380, Pix_381, Pix_382, Pix_383, Pix_384, Pix_385, Pix_386, Pix_387, Pix_388, Pix_389, Pix_390, Pix_391, Pix_392, Pix_393, Pix_394, Pix_395, Pix_396, Pix_397, Pix_398, Pix_399, Pix_400, Pix_401, Pix_402, Pix_403, Pix_404, Pix_405, Pix_406, Pix_407, Pix_408, Pix_409, Pix_410, Pix_411, Pix_412, Pix_413, Pix_414, Pix_415, Pix_416, Pix_417, Pix_418, Pix_419, Pix_420, Pix_421, Pix_422, Pix_423, Pix_424, Pix_425, Pix_426, Pix_427, Pix_428, Pix_429, Pix_430, Pix_431, Pix_432, Pix_433, Pix_434, Pix_435, Pix_436, Pix_437, Pix_438, Pix_439, Pix_440, Pix_441, Pix_442, Pix_443, Pix_444, Pix_445, Pix_446, Pix_447, Pix_448, Pix_449, Pix_450, Pix_451, Pix_452, Pix_453, Pix_454, Pix_455, Pix_456, Pix_457, Pix_458, Pix_459, Pix_460, Pix_461, Pix_462, Pix_463, Pix_464, Pix_465, Pix_466, Pix_467, Pix_468, Pix_469, Pix_470, Pix_471, Pix_472, Pix_473, Pix_474, Pix_475, Pix_476, Pix_477, Pix_478, Pix_479, Pix_480, Pix_481, Pix_482, Pix_483, Pix_484, Pix_485, Pix_486, Pix_487, Pix_488, Pix_489, Pix_490, Pix_491, Pix_492, Pix_493, Pix_494, Pix_495, Pix_496, Pix_497, Pix_498, Pix_499, Pix_500, Pix_501, Pix_502, Pix_503, Pix_504, Pix_505, Pix_506, Pix_507, Pix_508, Pix_509, Pix_510, Pix_511, Pix_512, Pix_513, Pix_514, Pix_515, Pix_516, Pix_517, Pix_518, Pix_519, Pix_520, Pix_521, Pix_522, Pix_523, Pix_524, Pix_525, Pix_526, Pix_527, Pix_528, Pix_529, Pix_530, Pix_531, Pix_532, Pix_533, Pix_534, Pix_535, Pix_536, Pix_537, Pix_538, Pix_539, Pix_540, Pix_541, Pix_542, Pix_543, Pix_544, Pix_545, Pix_546, Pix_547, Pix_548, Pix_549, Pix_550, Pix_551, Pix_552, Pix_553, Pix_554, Pix_555, Pix_556, Pix_557, Pix_558, Pix_559, Pix_560, Pix_561, Pix_562, Pix_563, Pix_564, Pix_565, Pix_566, Pix_567, Pix_568, Pix_569, Pix_570, Pix_571, Pix_572, Pix_573, Pix_574, Pix_575, Pix_576, Pix_577, Pix_578, Pix_579, Pix_580, Pix_581, Pix_582, Pix_583, Pix_584, Pix_585, Pix_586, Pix_587, Pix_588, Pix_589, Pix_590, Pix_591, Pix_592, Pix_593, Pix_594, Pix_595, Pix_596, Pix_597, Pix_598, Pix_599, Pix_600, Pix_601, Pix_602, Pix_603, Pix_604, Pix_605, Pix_606, Pix_607, Pix_608, Pix_609, Pix_610, Pix_611, Pix_612, Pix_613, Pix_614, Pix_615, Pix_616, Pix_617, Pix_618, Pix_619, Pix_620, Pix_621, Pix_622, Pix_623, Pix_624, Pix_625, Pix_626, Pix_627, Pix_628, Pix_629, Pix_630, Pix_631, Pix_632, Pix_633, Pix_634, Pix_635, Pix_636, Pix_637, Pix_638, Pix_639, Pix_640, Pix_641, Pix_642, Pix_643, Pix_644, Pix_645, Pix_646, Pix_647, Pix_648, Pix_649, Pix_650, Pix_651, Pix_652, Pix_653, Pix_654, Pix_655, Pix_656, Pix_657, Pix_658, Pix_659, Pix_660, Pix_661, Pix_662, Pix_663, Pix_664, Pix_665, Pix_666, Pix_667, Pix_668, Pix_669, Pix_670, Pix_671, Pix_672, Pix_673, Pix_674, Pix_675, Pix_676, Pix_677, Pix_678, Pix_679, Pix_680, Pix_681, Pix_682, Pix_683, Pix_684, Pix_685, Pix_686, Pix_687, Pix_688, Pix_689, Pix_690, Pix_691, Pix_692, Pix_693, Pix_694, Pix_695, Pix_696, Pix_697, Pix_698, Pix_699, Pix_700, Pix_701, Pix_702, Pix_703, Pix_704, Pix_705, Pix_706, Pix_707, Pix_708, Pix_709, Pix_710, Pix_711, Pix_712, Pix_713, Pix_714, Pix_715, Pix_716, Pix_717, Pix_718, Pix_719, Pix_720, Pix_721, Pix_722, Pix_723, Pix_724, Pix_725, Pix_726, Pix_727, Pix_728, Pix_729, Pix_730, Pix_731, Pix_732, Pix_733, Pix_734, Pix_735, Pix_736, Pix_737, Pix_738, Pix_739, Pix_740, Pix_741, Pix_742, Pix_743, Pix_744, Pix_745, Pix_746, Pix_747, Pix_748, Pix_749, Pix_750, Pix_751, Pix_752, Pix_753, Pix_754, Pix_755, Pix_756, Pix_757, Pix_758, Pix_759, Pix_760, Pix_761, Pix_762, Pix_763, Pix_764, Pix_765, Pix_766, Pix_767, Pix_768, Pix_769, Pix_770, Pix_771, Pix_772, Pix_773, Pix_774, Pix_775, Pix_776, Pix_777, Pix_778, Pix_779, Pix_780, Pix_781, Pix_782, Pix_783,
	output reg [9:0] Pix_0_reg, Pix_1_reg, Pix_2_reg, Pix_3_reg, Pix_4_reg, Pix_5_reg, Pix_6_reg, Pix_7_reg, Pix_8_reg, Pix_9_reg, Pix_10_reg, Pix_11_reg, Pix_12_reg, Pix_13_reg, Pix_14_reg, Pix_15_reg, Pix_16_reg, Pix_17_reg, Pix_18_reg, Pix_19_reg, Pix_20_reg, Pix_21_reg, Pix_22_reg, Pix_23_reg, Pix_24_reg, Pix_25_reg, Pix_26_reg, Pix_27_reg, Pix_28_reg, Pix_29_reg, Pix_30_reg, Pix_31_reg, Pix_32_reg, Pix_33_reg, Pix_34_reg, Pix_35_reg, Pix_36_reg, Pix_37_reg, Pix_38_reg, Pix_39_reg, Pix_40_reg, Pix_41_reg, Pix_42_reg, Pix_43_reg, Pix_44_reg, Pix_45_reg, Pix_46_reg, Pix_47_reg, Pix_48_reg, Pix_49_reg, Pix_50_reg, Pix_51_reg, Pix_52_reg, Pix_53_reg, Pix_54_reg, Pix_55_reg, Pix_56_reg, Pix_57_reg, Pix_58_reg, Pix_59_reg, Pix_60_reg, Pix_61_reg, Pix_62_reg, Pix_63_reg, Pix_64_reg, Pix_65_reg, Pix_66_reg, Pix_67_reg, Pix_68_reg, Pix_69_reg, Pix_70_reg, Pix_71_reg, Pix_72_reg, Pix_73_reg, Pix_74_reg, Pix_75_reg, Pix_76_reg, Pix_77_reg, Pix_78_reg, Pix_79_reg, Pix_80_reg, Pix_81_reg, Pix_82_reg, Pix_83_reg, Pix_84_reg, Pix_85_reg, Pix_86_reg, Pix_87_reg, Pix_88_reg, Pix_89_reg, Pix_90_reg, Pix_91_reg, Pix_92_reg, Pix_93_reg, Pix_94_reg, Pix_95_reg, Pix_96_reg, Pix_97_reg, Pix_98_reg, Pix_99_reg, Pix_100_reg, Pix_101_reg, Pix_102_reg, Pix_103_reg, Pix_104_reg, Pix_105_reg, Pix_106_reg, Pix_107_reg, Pix_108_reg, Pix_109_reg, Pix_110_reg, Pix_111_reg, Pix_112_reg, Pix_113_reg, Pix_114_reg, Pix_115_reg, Pix_116_reg, Pix_117_reg, Pix_118_reg, Pix_119_reg, Pix_120_reg, Pix_121_reg, Pix_122_reg, Pix_123_reg, Pix_124_reg, Pix_125_reg, Pix_126_reg, Pix_127_reg, Pix_128_reg, Pix_129_reg, Pix_130_reg, Pix_131_reg, Pix_132_reg, Pix_133_reg, Pix_134_reg, Pix_135_reg, Pix_136_reg, Pix_137_reg, Pix_138_reg, Pix_139_reg, Pix_140_reg, Pix_141_reg, Pix_142_reg, Pix_143_reg, Pix_144_reg, Pix_145_reg, Pix_146_reg, Pix_147_reg, Pix_148_reg, Pix_149_reg, Pix_150_reg, Pix_151_reg, Pix_152_reg, Pix_153_reg, Pix_154_reg, Pix_155_reg, Pix_156_reg, Pix_157_reg, Pix_158_reg, Pix_159_reg, Pix_160_reg, Pix_161_reg, Pix_162_reg, Pix_163_reg, Pix_164_reg, Pix_165_reg, Pix_166_reg, Pix_167_reg, Pix_168_reg, Pix_169_reg, Pix_170_reg, Pix_171_reg, Pix_172_reg, Pix_173_reg, Pix_174_reg, Pix_175_reg, Pix_176_reg, Pix_177_reg, Pix_178_reg, Pix_179_reg, Pix_180_reg, Pix_181_reg, Pix_182_reg, Pix_183_reg, Pix_184_reg, Pix_185_reg, Pix_186_reg, Pix_187_reg, Pix_188_reg, Pix_189_reg, Pix_190_reg, Pix_191_reg, Pix_192_reg, Pix_193_reg, Pix_194_reg, Pix_195_reg, Pix_196_reg, Pix_197_reg, Pix_198_reg, Pix_199_reg, Pix_200_reg, Pix_201_reg, Pix_202_reg, Pix_203_reg, Pix_204_reg, Pix_205_reg, Pix_206_reg, Pix_207_reg, Pix_208_reg, Pix_209_reg, Pix_210_reg, Pix_211_reg, Pix_212_reg, Pix_213_reg, Pix_214_reg, Pix_215_reg, Pix_216_reg, Pix_217_reg, Pix_218_reg, Pix_219_reg, Pix_220_reg, Pix_221_reg, Pix_222_reg, Pix_223_reg, Pix_224_reg, Pix_225_reg, Pix_226_reg, Pix_227_reg, Pix_228_reg, Pix_229_reg, Pix_230_reg, Pix_231_reg, Pix_232_reg, Pix_233_reg, Pix_234_reg, Pix_235_reg, Pix_236_reg, Pix_237_reg, Pix_238_reg, Pix_239_reg, Pix_240_reg, Pix_241_reg, Pix_242_reg, Pix_243_reg, Pix_244_reg, Pix_245_reg, Pix_246_reg, Pix_247_reg, Pix_248_reg, Pix_249_reg, Pix_250_reg, Pix_251_reg, Pix_252_reg, Pix_253_reg, Pix_254_reg, Pix_255_reg, Pix_256_reg, Pix_257_reg, Pix_258_reg, Pix_259_reg, Pix_260_reg, Pix_261_reg, Pix_262_reg, Pix_263_reg, Pix_264_reg, Pix_265_reg, Pix_266_reg, Pix_267_reg, Pix_268_reg, Pix_269_reg, Pix_270_reg, Pix_271_reg, Pix_272_reg, Pix_273_reg, Pix_274_reg, Pix_275_reg, Pix_276_reg, Pix_277_reg, Pix_278_reg, Pix_279_reg, Pix_280_reg, Pix_281_reg, Pix_282_reg, Pix_283_reg, Pix_284_reg, Pix_285_reg, Pix_286_reg, Pix_287_reg, Pix_288_reg, Pix_289_reg, Pix_290_reg, Pix_291_reg, Pix_292_reg, Pix_293_reg, Pix_294_reg, Pix_295_reg, Pix_296_reg, Pix_297_reg, Pix_298_reg, Pix_299_reg, Pix_300_reg, Pix_301_reg, Pix_302_reg, Pix_303_reg, Pix_304_reg, Pix_305_reg, Pix_306_reg, Pix_307_reg, Pix_308_reg, Pix_309_reg, Pix_310_reg, Pix_311_reg, Pix_312_reg, Pix_313_reg, Pix_314_reg, Pix_315_reg, Pix_316_reg, Pix_317_reg, Pix_318_reg, Pix_319_reg, Pix_320_reg, Pix_321_reg, Pix_322_reg, Pix_323_reg, Pix_324_reg, Pix_325_reg, Pix_326_reg, Pix_327_reg, Pix_328_reg, Pix_329_reg, Pix_330_reg, Pix_331_reg, Pix_332_reg, Pix_333_reg, Pix_334_reg, Pix_335_reg, Pix_336_reg, Pix_337_reg, Pix_338_reg, Pix_339_reg, Pix_340_reg, Pix_341_reg, Pix_342_reg, Pix_343_reg, Pix_344_reg, Pix_345_reg, Pix_346_reg, Pix_347_reg, Pix_348_reg, Pix_349_reg, Pix_350_reg, Pix_351_reg, Pix_352_reg, Pix_353_reg, Pix_354_reg, Pix_355_reg, Pix_356_reg, Pix_357_reg, Pix_358_reg, Pix_359_reg, Pix_360_reg, Pix_361_reg, Pix_362_reg, Pix_363_reg, Pix_364_reg, Pix_365_reg, Pix_366_reg, Pix_367_reg, Pix_368_reg, Pix_369_reg, Pix_370_reg, Pix_371_reg, Pix_372_reg, Pix_373_reg, Pix_374_reg, Pix_375_reg, Pix_376_reg, Pix_377_reg, Pix_378_reg, Pix_379_reg, Pix_380_reg, Pix_381_reg, Pix_382_reg, Pix_383_reg, Pix_384_reg, Pix_385_reg, Pix_386_reg, Pix_387_reg, Pix_388_reg, Pix_389_reg, Pix_390_reg, Pix_391_reg, Pix_392_reg, Pix_393_reg, Pix_394_reg, Pix_395_reg, Pix_396_reg, Pix_397_reg, Pix_398_reg, Pix_399_reg, Pix_400_reg, Pix_401_reg, Pix_402_reg, Pix_403_reg, Pix_404_reg, Pix_405_reg, Pix_406_reg, Pix_407_reg, Pix_408_reg, Pix_409_reg, Pix_410_reg, Pix_411_reg, Pix_412_reg, Pix_413_reg, Pix_414_reg, Pix_415_reg, Pix_416_reg, Pix_417_reg, Pix_418_reg, Pix_419_reg, Pix_420_reg, Pix_421_reg, Pix_422_reg, Pix_423_reg, Pix_424_reg, Pix_425_reg, Pix_426_reg, Pix_427_reg, Pix_428_reg, Pix_429_reg, Pix_430_reg, Pix_431_reg, Pix_432_reg, Pix_433_reg, Pix_434_reg, Pix_435_reg, Pix_436_reg, Pix_437_reg, Pix_438_reg, Pix_439_reg, Pix_440_reg, Pix_441_reg, Pix_442_reg, Pix_443_reg, Pix_444_reg, Pix_445_reg, Pix_446_reg, Pix_447_reg, Pix_448_reg, Pix_449_reg, Pix_450_reg, Pix_451_reg, Pix_452_reg, Pix_453_reg, Pix_454_reg, Pix_455_reg, Pix_456_reg, Pix_457_reg, Pix_458_reg, Pix_459_reg, Pix_460_reg, Pix_461_reg, Pix_462_reg, Pix_463_reg, Pix_464_reg, Pix_465_reg, Pix_466_reg, Pix_467_reg, Pix_468_reg, Pix_469_reg, Pix_470_reg, Pix_471_reg, Pix_472_reg, Pix_473_reg, Pix_474_reg, Pix_475_reg, Pix_476_reg, Pix_477_reg, Pix_478_reg, Pix_479_reg, Pix_480_reg, Pix_481_reg, Pix_482_reg, Pix_483_reg, Pix_484_reg, Pix_485_reg, Pix_486_reg, Pix_487_reg, Pix_488_reg, Pix_489_reg, Pix_490_reg, Pix_491_reg, Pix_492_reg, Pix_493_reg, Pix_494_reg, Pix_495_reg, Pix_496_reg, Pix_497_reg, Pix_498_reg, Pix_499_reg, Pix_500_reg, Pix_501_reg, Pix_502_reg, Pix_503_reg, Pix_504_reg, Pix_505_reg, Pix_506_reg, Pix_507_reg, Pix_508_reg, Pix_509_reg, Pix_510_reg, Pix_511_reg, Pix_512_reg, Pix_513_reg, Pix_514_reg, Pix_515_reg, Pix_516_reg, Pix_517_reg, Pix_518_reg, Pix_519_reg, Pix_520_reg, Pix_521_reg, Pix_522_reg, Pix_523_reg, Pix_524_reg, Pix_525_reg, Pix_526_reg, Pix_527_reg, Pix_528_reg, Pix_529_reg, Pix_530_reg, Pix_531_reg, Pix_532_reg, Pix_533_reg, Pix_534_reg, Pix_535_reg, Pix_536_reg, Pix_537_reg, Pix_538_reg, Pix_539_reg, Pix_540_reg, Pix_541_reg, Pix_542_reg, Pix_543_reg, Pix_544_reg, Pix_545_reg, Pix_546_reg, Pix_547_reg, Pix_548_reg, Pix_549_reg, Pix_550_reg, Pix_551_reg, Pix_552_reg, Pix_553_reg, Pix_554_reg, Pix_555_reg, Pix_556_reg, Pix_557_reg, Pix_558_reg, Pix_559_reg, Pix_560_reg, Pix_561_reg, Pix_562_reg, Pix_563_reg, Pix_564_reg, Pix_565_reg, Pix_566_reg, Pix_567_reg, Pix_568_reg, Pix_569_reg, Pix_570_reg, Pix_571_reg, Pix_572_reg, Pix_573_reg, Pix_574_reg, Pix_575_reg, Pix_576_reg, Pix_577_reg, Pix_578_reg, Pix_579_reg, Pix_580_reg, Pix_581_reg, Pix_582_reg, Pix_583_reg, Pix_584_reg, Pix_585_reg, Pix_586_reg, Pix_587_reg, Pix_588_reg, Pix_589_reg, Pix_590_reg, Pix_591_reg, Pix_592_reg, Pix_593_reg, Pix_594_reg, Pix_595_reg, Pix_596_reg, Pix_597_reg, Pix_598_reg, Pix_599_reg, Pix_600_reg, Pix_601_reg, Pix_602_reg, Pix_603_reg, Pix_604_reg, Pix_605_reg, Pix_606_reg, Pix_607_reg, Pix_608_reg, Pix_609_reg, Pix_610_reg, Pix_611_reg, Pix_612_reg, Pix_613_reg, Pix_614_reg, Pix_615_reg, Pix_616_reg, Pix_617_reg, Pix_618_reg, Pix_619_reg, Pix_620_reg, Pix_621_reg, Pix_622_reg, Pix_623_reg, Pix_624_reg, Pix_625_reg, Pix_626_reg, Pix_627_reg, Pix_628_reg, Pix_629_reg, Pix_630_reg, Pix_631_reg, Pix_632_reg, Pix_633_reg, Pix_634_reg, Pix_635_reg, Pix_636_reg, Pix_637_reg, Pix_638_reg, Pix_639_reg, Pix_640_reg, Pix_641_reg, Pix_642_reg, Pix_643_reg, Pix_644_reg, Pix_645_reg, Pix_646_reg, Pix_647_reg, Pix_648_reg, Pix_649_reg, Pix_650_reg, Pix_651_reg, Pix_652_reg, Pix_653_reg, Pix_654_reg, Pix_655_reg, Pix_656_reg, Pix_657_reg, Pix_658_reg, Pix_659_reg, Pix_660_reg, Pix_661_reg, Pix_662_reg, Pix_663_reg, Pix_664_reg, Pix_665_reg, Pix_666_reg, Pix_667_reg, Pix_668_reg, Pix_669_reg, Pix_670_reg, Pix_671_reg, Pix_672_reg, Pix_673_reg, Pix_674_reg, Pix_675_reg, Pix_676_reg, Pix_677_reg, Pix_678_reg, Pix_679_reg, Pix_680_reg, Pix_681_reg, Pix_682_reg, Pix_683_reg, Pix_684_reg, Pix_685_reg, Pix_686_reg, Pix_687_reg, Pix_688_reg, Pix_689_reg, Pix_690_reg, Pix_691_reg, Pix_692_reg, Pix_693_reg, Pix_694_reg, Pix_695_reg, Pix_696_reg, Pix_697_reg, Pix_698_reg, Pix_699_reg, Pix_700_reg, Pix_701_reg, Pix_702_reg, Pix_703_reg, Pix_704_reg, Pix_705_reg, Pix_706_reg, Pix_707_reg, Pix_708_reg, Pix_709_reg, Pix_710_reg, Pix_711_reg, Pix_712_reg, Pix_713_reg, Pix_714_reg, Pix_715_reg, Pix_716_reg, Pix_717_reg, Pix_718_reg, Pix_719_reg, Pix_720_reg, Pix_721_reg, Pix_722_reg, Pix_723_reg, Pix_724_reg, Pix_725_reg, Pix_726_reg, Pix_727_reg, Pix_728_reg, Pix_729_reg, Pix_730_reg, Pix_731_reg, Pix_732_reg, Pix_733_reg, Pix_734_reg, Pix_735_reg, Pix_736_reg, Pix_737_reg, Pix_738_reg, Pix_739_reg, Pix_740_reg, Pix_741_reg, Pix_742_reg, Pix_743_reg, Pix_744_reg, Pix_745_reg, Pix_746_reg, Pix_747_reg, Pix_748_reg, Pix_749_reg, Pix_750_reg, Pix_751_reg, Pix_752_reg, Pix_753_reg, Pix_754_reg, Pix_755_reg, Pix_756_reg, Pix_757_reg, Pix_758_reg, Pix_759_reg, Pix_760_reg, Pix_761_reg, Pix_762_reg, Pix_763_reg, Pix_764_reg, Pix_765_reg, Pix_766_reg, Pix_767_reg, Pix_768_reg, Pix_769_reg, Pix_770_reg, Pix_771_reg, Pix_772_reg, Pix_773_reg, Pix_774_reg, Pix_775_reg, Pix_776_reg, Pix_777_reg, Pix_778_reg, Pix_779_reg, Pix_780_reg, Pix_781_reg, Pix_782_reg, Pix_783_reg );
	
	always @ (posedge clk) begin
		if (enable) begin
			 Pix_0_reg <= Pix_0;
			 Pix_1_reg <= Pix_1;
			 Pix_2_reg <= Pix_2;
			 Pix_3_reg <= Pix_3;
			 Pix_4_reg <= Pix_4;
			 Pix_5_reg <= Pix_5;
			 Pix_6_reg <= Pix_6;
			 Pix_7_reg <= Pix_7;
			 Pix_8_reg <= Pix_8;
			 Pix_9_reg <= Pix_9;
			 Pix_10_reg <= Pix_10;
			 Pix_11_reg <= Pix_11;
			 Pix_12_reg <= Pix_12;
			 Pix_13_reg <= Pix_13;
			 Pix_14_reg <= Pix_14;
			 Pix_15_reg <= Pix_15;
			 Pix_16_reg <= Pix_16;
			 Pix_17_reg <= Pix_17;
			 Pix_18_reg <= Pix_18;
			 Pix_19_reg <= Pix_19;
			 Pix_20_reg <= Pix_20;
			 Pix_21_reg <= Pix_21;
			 Pix_22_reg <= Pix_22;
			 Pix_23_reg <= Pix_23;
			 Pix_24_reg <= Pix_24;
			 Pix_25_reg <= Pix_25;
			 Pix_26_reg <= Pix_26;
			 Pix_27_reg <= Pix_27;
			 Pix_28_reg <= Pix_28;
			 Pix_29_reg <= Pix_29;
			 Pix_30_reg <= Pix_30;
			 Pix_31_reg <= Pix_31;
			 Pix_32_reg <= Pix_32;
			 Pix_33_reg <= Pix_33;
			 Pix_34_reg <= Pix_34;
			 Pix_35_reg <= Pix_35;
			 Pix_36_reg <= Pix_36;
			 Pix_37_reg <= Pix_37;
			 Pix_38_reg <= Pix_38;
			 Pix_39_reg <= Pix_39;
			 Pix_40_reg <= Pix_40;
			 Pix_41_reg <= Pix_41;
			 Pix_42_reg <= Pix_42;
			 Pix_43_reg <= Pix_43;
			 Pix_44_reg <= Pix_44;
			 Pix_45_reg <= Pix_45;
			 Pix_46_reg <= Pix_46;
			 Pix_47_reg <= Pix_47;
			 Pix_48_reg <= Pix_48;
			 Pix_49_reg <= Pix_49;
			 Pix_50_reg <= Pix_50;
			 Pix_51_reg <= Pix_51;
			 Pix_52_reg <= Pix_52;
			 Pix_53_reg <= Pix_53;
			 Pix_54_reg <= Pix_54;
			 Pix_55_reg <= Pix_55;
			 Pix_56_reg <= Pix_56;
			 Pix_57_reg <= Pix_57;
			 Pix_58_reg <= Pix_58;
			 Pix_59_reg <= Pix_59;
			 Pix_60_reg <= Pix_60;
			 Pix_61_reg <= Pix_61;
			 Pix_62_reg <= Pix_62;
			 Pix_63_reg <= Pix_63;
			 Pix_64_reg <= Pix_64;
			 Pix_65_reg <= Pix_65;
			 Pix_66_reg <= Pix_66;
			 Pix_67_reg <= Pix_67;
			 Pix_68_reg <= Pix_68;
			 Pix_69_reg <= Pix_69;
			 Pix_70_reg <= Pix_70;
			 Pix_71_reg <= Pix_71;
			 Pix_72_reg <= Pix_72;
			 Pix_73_reg <= Pix_73;
			 Pix_74_reg <= Pix_74;
			 Pix_75_reg <= Pix_75;
			 Pix_76_reg <= Pix_76;
			 Pix_77_reg <= Pix_77;
			 Pix_78_reg <= Pix_78;
			 Pix_79_reg <= Pix_79;
			 Pix_80_reg <= Pix_80;
			 Pix_81_reg <= Pix_81;
			 Pix_82_reg <= Pix_82;
			 Pix_83_reg <= Pix_83;
			 Pix_84_reg <= Pix_84;
			 Pix_85_reg <= Pix_85;
			 Pix_86_reg <= Pix_86;
			 Pix_87_reg <= Pix_87;
			 Pix_88_reg <= Pix_88;
			 Pix_89_reg <= Pix_89;
			 Pix_90_reg <= Pix_90;
			 Pix_91_reg <= Pix_91;
			 Pix_92_reg <= Pix_92;
			 Pix_93_reg <= Pix_93;
			 Pix_94_reg <= Pix_94;
			 Pix_95_reg <= Pix_95;
			 Pix_96_reg <= Pix_96;
			 Pix_97_reg <= Pix_97;
			 Pix_98_reg <= Pix_98;
			 Pix_99_reg <= Pix_99;
			 Pix_100_reg <= Pix_100;
			 Pix_101_reg <= Pix_101;
			 Pix_102_reg <= Pix_102;
			 Pix_103_reg <= Pix_103;
			 Pix_104_reg <= Pix_104;
			 Pix_105_reg <= Pix_105;
			 Pix_106_reg <= Pix_106;
			 Pix_107_reg <= Pix_107;
			 Pix_108_reg <= Pix_108;
			 Pix_109_reg <= Pix_109;
			 Pix_110_reg <= Pix_110;
			 Pix_111_reg <= Pix_111;
			 Pix_112_reg <= Pix_112;
			 Pix_113_reg <= Pix_113;
			 Pix_114_reg <= Pix_114;
			 Pix_115_reg <= Pix_115;
			 Pix_116_reg <= Pix_116;
			 Pix_117_reg <= Pix_117;
			 Pix_118_reg <= Pix_118;
			 Pix_119_reg <= Pix_119;
			 Pix_120_reg <= Pix_120;
			 Pix_121_reg <= Pix_121;
			 Pix_122_reg <= Pix_122;
			 Pix_123_reg <= Pix_123;
			 Pix_124_reg <= Pix_124;
			 Pix_125_reg <= Pix_125;
			 Pix_126_reg <= Pix_126;
			 Pix_127_reg <= Pix_127;
			 Pix_128_reg <= Pix_128;
			 Pix_129_reg <= Pix_129;
			 Pix_130_reg <= Pix_130;
			 Pix_131_reg <= Pix_131;
			 Pix_132_reg <= Pix_132;
			 Pix_133_reg <= Pix_133;
			 Pix_134_reg <= Pix_134;
			 Pix_135_reg <= Pix_135;
			 Pix_136_reg <= Pix_136;
			 Pix_137_reg <= Pix_137;
			 Pix_138_reg <= Pix_138;
			 Pix_139_reg <= Pix_139;
			 Pix_140_reg <= Pix_140;
			 Pix_141_reg <= Pix_141;
			 Pix_142_reg <= Pix_142;
			 Pix_143_reg <= Pix_143;
			 Pix_144_reg <= Pix_144;
			 Pix_145_reg <= Pix_145;
			 Pix_146_reg <= Pix_146;
			 Pix_147_reg <= Pix_147;
			 Pix_148_reg <= Pix_148;
			 Pix_149_reg <= Pix_149;
			 Pix_150_reg <= Pix_150;
			 Pix_151_reg <= Pix_151;
			 Pix_152_reg <= Pix_152;
			 Pix_153_reg <= Pix_153;
			 Pix_154_reg <= Pix_154;
			 Pix_155_reg <= Pix_155;
			 Pix_156_reg <= Pix_156;
			 Pix_157_reg <= Pix_157;
			 Pix_158_reg <= Pix_158;
			 Pix_159_reg <= Pix_159;
			 Pix_160_reg <= Pix_160;
			 Pix_161_reg <= Pix_161;
			 Pix_162_reg <= Pix_162;
			 Pix_163_reg <= Pix_163;
			 Pix_164_reg <= Pix_164;
			 Pix_165_reg <= Pix_165;
			 Pix_166_reg <= Pix_166;
			 Pix_167_reg <= Pix_167;
			 Pix_168_reg <= Pix_168;
			 Pix_169_reg <= Pix_169;
			 Pix_170_reg <= Pix_170;
			 Pix_171_reg <= Pix_171;
			 Pix_172_reg <= Pix_172;
			 Pix_173_reg <= Pix_173;
			 Pix_174_reg <= Pix_174;
			 Pix_175_reg <= Pix_175;
			 Pix_176_reg <= Pix_176;
			 Pix_177_reg <= Pix_177;
			 Pix_178_reg <= Pix_178;
			 Pix_179_reg <= Pix_179;
			 Pix_180_reg <= Pix_180;
			 Pix_181_reg <= Pix_181;
			 Pix_182_reg <= Pix_182;
			 Pix_183_reg <= Pix_183;
			 Pix_184_reg <= Pix_184;
			 Pix_185_reg <= Pix_185;
			 Pix_186_reg <= Pix_186;
			 Pix_187_reg <= Pix_187;
			 Pix_188_reg <= Pix_188;
			 Pix_189_reg <= Pix_189;
			 Pix_190_reg <= Pix_190;
			 Pix_191_reg <= Pix_191;
			 Pix_192_reg <= Pix_192;
			 Pix_193_reg <= Pix_193;
			 Pix_194_reg <= Pix_194;
			 Pix_195_reg <= Pix_195;
			 Pix_196_reg <= Pix_196;
			 Pix_197_reg <= Pix_197;
			 Pix_198_reg <= Pix_198;
			 Pix_199_reg <= Pix_199;
			 Pix_200_reg <= Pix_200;
			 Pix_201_reg <= Pix_201;
			 Pix_202_reg <= Pix_202;
			 Pix_203_reg <= Pix_203;
			 Pix_204_reg <= Pix_204;
			 Pix_205_reg <= Pix_205;
			 Pix_206_reg <= Pix_206;
			 Pix_207_reg <= Pix_207;
			 Pix_208_reg <= Pix_208;
			 Pix_209_reg <= Pix_209;
			 Pix_210_reg <= Pix_210;
			 Pix_211_reg <= Pix_211;
			 Pix_212_reg <= Pix_212;
			 Pix_213_reg <= Pix_213;
			 Pix_214_reg <= Pix_214;
			 Pix_215_reg <= Pix_215;
			 Pix_216_reg <= Pix_216;
			 Pix_217_reg <= Pix_217;
			 Pix_218_reg <= Pix_218;
			 Pix_219_reg <= Pix_219;
			 Pix_220_reg <= Pix_220;
			 Pix_221_reg <= Pix_221;
			 Pix_222_reg <= Pix_222;
			 Pix_223_reg <= Pix_223;
			 Pix_224_reg <= Pix_224;
			 Pix_225_reg <= Pix_225;
			 Pix_226_reg <= Pix_226;
			 Pix_227_reg <= Pix_227;
			 Pix_228_reg <= Pix_228;
			 Pix_229_reg <= Pix_229;
			 Pix_230_reg <= Pix_230;
			 Pix_231_reg <= Pix_231;
			 Pix_232_reg <= Pix_232;
			 Pix_233_reg <= Pix_233;
			 Pix_234_reg <= Pix_234;
			 Pix_235_reg <= Pix_235;
			 Pix_236_reg <= Pix_236;
			 Pix_237_reg <= Pix_237;
			 Pix_238_reg <= Pix_238;
			 Pix_239_reg <= Pix_239;
			 Pix_240_reg <= Pix_240;
			 Pix_241_reg <= Pix_241;
			 Pix_242_reg <= Pix_242;
			 Pix_243_reg <= Pix_243;
			 Pix_244_reg <= Pix_244;
			 Pix_245_reg <= Pix_245;
			 Pix_246_reg <= Pix_246;
			 Pix_247_reg <= Pix_247;
			 Pix_248_reg <= Pix_248;
			 Pix_249_reg <= Pix_249;
			 Pix_250_reg <= Pix_250;
			 Pix_251_reg <= Pix_251;
			 Pix_252_reg <= Pix_252;
			 Pix_253_reg <= Pix_253;
			 Pix_254_reg <= Pix_254;
			 Pix_255_reg <= Pix_255;
			 Pix_256_reg <= Pix_256;
			 Pix_257_reg <= Pix_257;
			 Pix_258_reg <= Pix_258;
			 Pix_259_reg <= Pix_259;
			 Pix_260_reg <= Pix_260;
			 Pix_261_reg <= Pix_261;
			 Pix_262_reg <= Pix_262;
			 Pix_263_reg <= Pix_263;
			 Pix_264_reg <= Pix_264;
			 Pix_265_reg <= Pix_265;
			 Pix_266_reg <= Pix_266;
			 Pix_267_reg <= Pix_267;
			 Pix_268_reg <= Pix_268;
			 Pix_269_reg <= Pix_269;
			 Pix_270_reg <= Pix_270;
			 Pix_271_reg <= Pix_271;
			 Pix_272_reg <= Pix_272;
			 Pix_273_reg <= Pix_273;
			 Pix_274_reg <= Pix_274;
			 Pix_275_reg <= Pix_275;
			 Pix_276_reg <= Pix_276;
			 Pix_277_reg <= Pix_277;
			 Pix_278_reg <= Pix_278;
			 Pix_279_reg <= Pix_279;
			 Pix_280_reg <= Pix_280;
			 Pix_281_reg <= Pix_281;
			 Pix_282_reg <= Pix_282;
			 Pix_283_reg <= Pix_283;
			 Pix_284_reg <= Pix_284;
			 Pix_285_reg <= Pix_285;
			 Pix_286_reg <= Pix_286;
			 Pix_287_reg <= Pix_287;
			 Pix_288_reg <= Pix_288;
			 Pix_289_reg <= Pix_289;
			 Pix_290_reg <= Pix_290;
			 Pix_291_reg <= Pix_291;
			 Pix_292_reg <= Pix_292;
			 Pix_293_reg <= Pix_293;
			 Pix_294_reg <= Pix_294;
			 Pix_295_reg <= Pix_295;
			 Pix_296_reg <= Pix_296;
			 Pix_297_reg <= Pix_297;
			 Pix_298_reg <= Pix_298;
			 Pix_299_reg <= Pix_299;
			 Pix_300_reg <= Pix_300;
			 Pix_301_reg <= Pix_301;
			 Pix_302_reg <= Pix_302;
			 Pix_303_reg <= Pix_303;
			 Pix_304_reg <= Pix_304;
			 Pix_305_reg <= Pix_305;
			 Pix_306_reg <= Pix_306;
			 Pix_307_reg <= Pix_307;
			 Pix_308_reg <= Pix_308;
			 Pix_309_reg <= Pix_309;
			 Pix_310_reg <= Pix_310;
			 Pix_311_reg <= Pix_311;
			 Pix_312_reg <= Pix_312;
			 Pix_313_reg <= Pix_313;
			 Pix_314_reg <= Pix_314;
			 Pix_315_reg <= Pix_315;
			 Pix_316_reg <= Pix_316;
			 Pix_317_reg <= Pix_317;
			 Pix_318_reg <= Pix_318;
			 Pix_319_reg <= Pix_319;
			 Pix_320_reg <= Pix_320;
			 Pix_321_reg <= Pix_321;
			 Pix_322_reg <= Pix_322;
			 Pix_323_reg <= Pix_323;
			 Pix_324_reg <= Pix_324;
			 Pix_325_reg <= Pix_325;
			 Pix_326_reg <= Pix_326;
			 Pix_327_reg <= Pix_327;
			 Pix_328_reg <= Pix_328;
			 Pix_329_reg <= Pix_329;
			 Pix_330_reg <= Pix_330;
			 Pix_331_reg <= Pix_331;
			 Pix_332_reg <= Pix_332;
			 Pix_333_reg <= Pix_333;
			 Pix_334_reg <= Pix_334;
			 Pix_335_reg <= Pix_335;
			 Pix_336_reg <= Pix_336;
			 Pix_337_reg <= Pix_337;
			 Pix_338_reg <= Pix_338;
			 Pix_339_reg <= Pix_339;
			 Pix_340_reg <= Pix_340;
			 Pix_341_reg <= Pix_341;
			 Pix_342_reg <= Pix_342;
			 Pix_343_reg <= Pix_343;
			 Pix_344_reg <= Pix_344;
			 Pix_345_reg <= Pix_345;
			 Pix_346_reg <= Pix_346;
			 Pix_347_reg <= Pix_347;
			 Pix_348_reg <= Pix_348;
			 Pix_349_reg <= Pix_349;
			 Pix_350_reg <= Pix_350;
			 Pix_351_reg <= Pix_351;
			 Pix_352_reg <= Pix_352;
			 Pix_353_reg <= Pix_353;
			 Pix_354_reg <= Pix_354;
			 Pix_355_reg <= Pix_355;
			 Pix_356_reg <= Pix_356;
			 Pix_357_reg <= Pix_357;
			 Pix_358_reg <= Pix_358;
			 Pix_359_reg <= Pix_359;
			 Pix_360_reg <= Pix_360;
			 Pix_361_reg <= Pix_361;
			 Pix_362_reg <= Pix_362;
			 Pix_363_reg <= Pix_363;
			 Pix_364_reg <= Pix_364;
			 Pix_365_reg <= Pix_365;
			 Pix_366_reg <= Pix_366;
			 Pix_367_reg <= Pix_367;
			 Pix_368_reg <= Pix_368;
			 Pix_369_reg <= Pix_369;
			 Pix_370_reg <= Pix_370;
			 Pix_371_reg <= Pix_371;
			 Pix_372_reg <= Pix_372;
			 Pix_373_reg <= Pix_373;
			 Pix_374_reg <= Pix_374;
			 Pix_375_reg <= Pix_375;
			 Pix_376_reg <= Pix_376;
			 Pix_377_reg <= Pix_377;
			 Pix_378_reg <= Pix_378;
			 Pix_379_reg <= Pix_379;
			 Pix_380_reg <= Pix_380;
			 Pix_381_reg <= Pix_381;
			 Pix_382_reg <= Pix_382;
			 Pix_383_reg <= Pix_383;
			 Pix_384_reg <= Pix_384;
			 Pix_385_reg <= Pix_385;
			 Pix_386_reg <= Pix_386;
			 Pix_387_reg <= Pix_387;
			 Pix_388_reg <= Pix_388;
			 Pix_389_reg <= Pix_389;
			 Pix_390_reg <= Pix_390;
			 Pix_391_reg <= Pix_391;
			 Pix_392_reg <= Pix_392;
			 Pix_393_reg <= Pix_393;
			 Pix_394_reg <= Pix_394;
			 Pix_395_reg <= Pix_395;
			 Pix_396_reg <= Pix_396;
			 Pix_397_reg <= Pix_397;
			 Pix_398_reg <= Pix_398;
			 Pix_399_reg <= Pix_399;
			 Pix_400_reg <= Pix_400;
			 Pix_401_reg <= Pix_401;
			 Pix_402_reg <= Pix_402;
			 Pix_403_reg <= Pix_403;
			 Pix_404_reg <= Pix_404;
			 Pix_405_reg <= Pix_405;
			 Pix_406_reg <= Pix_406;
			 Pix_407_reg <= Pix_407;
			 Pix_408_reg <= Pix_408;
			 Pix_409_reg <= Pix_409;
			 Pix_410_reg <= Pix_410;
			 Pix_411_reg <= Pix_411;
			 Pix_412_reg <= Pix_412;
			 Pix_413_reg <= Pix_413;
			 Pix_414_reg <= Pix_414;
			 Pix_415_reg <= Pix_415;
			 Pix_416_reg <= Pix_416;
			 Pix_417_reg <= Pix_417;
			 Pix_418_reg <= Pix_418;
			 Pix_419_reg <= Pix_419;
			 Pix_420_reg <= Pix_420;
			 Pix_421_reg <= Pix_421;
			 Pix_422_reg <= Pix_422;
			 Pix_423_reg <= Pix_423;
			 Pix_424_reg <= Pix_424;
			 Pix_425_reg <= Pix_425;
			 Pix_426_reg <= Pix_426;
			 Pix_427_reg <= Pix_427;
			 Pix_428_reg <= Pix_428;
			 Pix_429_reg <= Pix_429;
			 Pix_430_reg <= Pix_430;
			 Pix_431_reg <= Pix_431;
			 Pix_432_reg <= Pix_432;
			 Pix_433_reg <= Pix_433;
			 Pix_434_reg <= Pix_434;
			 Pix_435_reg <= Pix_435;
			 Pix_436_reg <= Pix_436;
			 Pix_437_reg <= Pix_437;
			 Pix_438_reg <= Pix_438;
			 Pix_439_reg <= Pix_439;
			 Pix_440_reg <= Pix_440;
			 Pix_441_reg <= Pix_441;
			 Pix_442_reg <= Pix_442;
			 Pix_443_reg <= Pix_443;
			 Pix_444_reg <= Pix_444;
			 Pix_445_reg <= Pix_445;
			 Pix_446_reg <= Pix_446;
			 Pix_447_reg <= Pix_447;
			 Pix_448_reg <= Pix_448;
			 Pix_449_reg <= Pix_449;
			 Pix_450_reg <= Pix_450;
			 Pix_451_reg <= Pix_451;
			 Pix_452_reg <= Pix_452;
			 Pix_453_reg <= Pix_453;
			 Pix_454_reg <= Pix_454;
			 Pix_455_reg <= Pix_455;
			 Pix_456_reg <= Pix_456;
			 Pix_457_reg <= Pix_457;
			 Pix_458_reg <= Pix_458;
			 Pix_459_reg <= Pix_459;
			 Pix_460_reg <= Pix_460;
			 Pix_461_reg <= Pix_461;
			 Pix_462_reg <= Pix_462;
			 Pix_463_reg <= Pix_463;
			 Pix_464_reg <= Pix_464;
			 Pix_465_reg <= Pix_465;
			 Pix_466_reg <= Pix_466;
			 Pix_467_reg <= Pix_467;
			 Pix_468_reg <= Pix_468;
			 Pix_469_reg <= Pix_469;
			 Pix_470_reg <= Pix_470;
			 Pix_471_reg <= Pix_471;
			 Pix_472_reg <= Pix_472;
			 Pix_473_reg <= Pix_473;
			 Pix_474_reg <= Pix_474;
			 Pix_475_reg <= Pix_475;
			 Pix_476_reg <= Pix_476;
			 Pix_477_reg <= Pix_477;
			 Pix_478_reg <= Pix_478;
			 Pix_479_reg <= Pix_479;
			 Pix_480_reg <= Pix_480;
			 Pix_481_reg <= Pix_481;
			 Pix_482_reg <= Pix_482;
			 Pix_483_reg <= Pix_483;
			 Pix_484_reg <= Pix_484;
			 Pix_485_reg <= Pix_485;
			 Pix_486_reg <= Pix_486;
			 Pix_487_reg <= Pix_487;
			 Pix_488_reg <= Pix_488;
			 Pix_489_reg <= Pix_489;
			 Pix_490_reg <= Pix_490;
			 Pix_491_reg <= Pix_491;
			 Pix_492_reg <= Pix_492;
			 Pix_493_reg <= Pix_493;
			 Pix_494_reg <= Pix_494;
			 Pix_495_reg <= Pix_495;
			 Pix_496_reg <= Pix_496;
			 Pix_497_reg <= Pix_497;
			 Pix_498_reg <= Pix_498;
			 Pix_499_reg <= Pix_499;
			 Pix_500_reg <= Pix_500;
			 Pix_501_reg <= Pix_501;
			 Pix_502_reg <= Pix_502;
			 Pix_503_reg <= Pix_503;
			 Pix_504_reg <= Pix_504;
			 Pix_505_reg <= Pix_505;
			 Pix_506_reg <= Pix_506;
			 Pix_507_reg <= Pix_507;
			 Pix_508_reg <= Pix_508;
			 Pix_509_reg <= Pix_509;
			 Pix_510_reg <= Pix_510;
			 Pix_511_reg <= Pix_511;
			 Pix_512_reg <= Pix_512;
			 Pix_513_reg <= Pix_513;
			 Pix_514_reg <= Pix_514;
			 Pix_515_reg <= Pix_515;
			 Pix_516_reg <= Pix_516;
			 Pix_517_reg <= Pix_517;
			 Pix_518_reg <= Pix_518;
			 Pix_519_reg <= Pix_519;
			 Pix_520_reg <= Pix_520;
			 Pix_521_reg <= Pix_521;
			 Pix_522_reg <= Pix_522;
			 Pix_523_reg <= Pix_523;
			 Pix_524_reg <= Pix_524;
			 Pix_525_reg <= Pix_525;
			 Pix_526_reg <= Pix_526;
			 Pix_527_reg <= Pix_527;
			 Pix_528_reg <= Pix_528;
			 Pix_529_reg <= Pix_529;
			 Pix_530_reg <= Pix_530;
			 Pix_531_reg <= Pix_531;
			 Pix_532_reg <= Pix_532;
			 Pix_533_reg <= Pix_533;
			 Pix_534_reg <= Pix_534;
			 Pix_535_reg <= Pix_535;
			 Pix_536_reg <= Pix_536;
			 Pix_537_reg <= Pix_537;
			 Pix_538_reg <= Pix_538;
			 Pix_539_reg <= Pix_539;
			 Pix_540_reg <= Pix_540;
			 Pix_541_reg <= Pix_541;
			 Pix_542_reg <= Pix_542;
			 Pix_543_reg <= Pix_543;
			 Pix_544_reg <= Pix_544;
			 Pix_545_reg <= Pix_545;
			 Pix_546_reg <= Pix_546;
			 Pix_547_reg <= Pix_547;
			 Pix_548_reg <= Pix_548;
			 Pix_549_reg <= Pix_549;
			 Pix_550_reg <= Pix_550;
			 Pix_551_reg <= Pix_551;
			 Pix_552_reg <= Pix_552;
			 Pix_553_reg <= Pix_553;
			 Pix_554_reg <= Pix_554;
			 Pix_555_reg <= Pix_555;
			 Pix_556_reg <= Pix_556;
			 Pix_557_reg <= Pix_557;
			 Pix_558_reg <= Pix_558;
			 Pix_559_reg <= Pix_559;
			 Pix_560_reg <= Pix_560;
			 Pix_561_reg <= Pix_561;
			 Pix_562_reg <= Pix_562;
			 Pix_563_reg <= Pix_563;
			 Pix_564_reg <= Pix_564;
			 Pix_565_reg <= Pix_565;
			 Pix_566_reg <= Pix_566;
			 Pix_567_reg <= Pix_567;
			 Pix_568_reg <= Pix_568;
			 Pix_569_reg <= Pix_569;
			 Pix_570_reg <= Pix_570;
			 Pix_571_reg <= Pix_571;
			 Pix_572_reg <= Pix_572;
			 Pix_573_reg <= Pix_573;
			 Pix_574_reg <= Pix_574;
			 Pix_575_reg <= Pix_575;
			 Pix_576_reg <= Pix_576;
			 Pix_577_reg <= Pix_577;
			 Pix_578_reg <= Pix_578;
			 Pix_579_reg <= Pix_579;
			 Pix_580_reg <= Pix_580;
			 Pix_581_reg <= Pix_581;
			 Pix_582_reg <= Pix_582;
			 Pix_583_reg <= Pix_583;
			 Pix_584_reg <= Pix_584;
			 Pix_585_reg <= Pix_585;
			 Pix_586_reg <= Pix_586;
			 Pix_587_reg <= Pix_587;
			 Pix_588_reg <= Pix_588;
			 Pix_589_reg <= Pix_589;
			 Pix_590_reg <= Pix_590;
			 Pix_591_reg <= Pix_591;
			 Pix_592_reg <= Pix_592;
			 Pix_593_reg <= Pix_593;
			 Pix_594_reg <= Pix_594;
			 Pix_595_reg <= Pix_595;
			 Pix_596_reg <= Pix_596;
			 Pix_597_reg <= Pix_597;
			 Pix_598_reg <= Pix_598;
			 Pix_599_reg <= Pix_599;
			 Pix_600_reg <= Pix_600;
			 Pix_601_reg <= Pix_601;
			 Pix_602_reg <= Pix_602;
			 Pix_603_reg <= Pix_603;
			 Pix_604_reg <= Pix_604;
			 Pix_605_reg <= Pix_605;
			 Pix_606_reg <= Pix_606;
			 Pix_607_reg <= Pix_607;
			 Pix_608_reg <= Pix_608;
			 Pix_609_reg <= Pix_609;
			 Pix_610_reg <= Pix_610;
			 Pix_611_reg <= Pix_611;
			 Pix_612_reg <= Pix_612;
			 Pix_613_reg <= Pix_613;
			 Pix_614_reg <= Pix_614;
			 Pix_615_reg <= Pix_615;
			 Pix_616_reg <= Pix_616;
			 Pix_617_reg <= Pix_617;
			 Pix_618_reg <= Pix_618;
			 Pix_619_reg <= Pix_619;
			 Pix_620_reg <= Pix_620;
			 Pix_621_reg <= Pix_621;
			 Pix_622_reg <= Pix_622;
			 Pix_623_reg <= Pix_623;
			 Pix_624_reg <= Pix_624;
			 Pix_625_reg <= Pix_625;
			 Pix_626_reg <= Pix_626;
			 Pix_627_reg <= Pix_627;
			 Pix_628_reg <= Pix_628;
			 Pix_629_reg <= Pix_629;
			 Pix_630_reg <= Pix_630;
			 Pix_631_reg <= Pix_631;
			 Pix_632_reg <= Pix_632;
			 Pix_633_reg <= Pix_633;
			 Pix_634_reg <= Pix_634;
			 Pix_635_reg <= Pix_635;
			 Pix_636_reg <= Pix_636;
			 Pix_637_reg <= Pix_637;
			 Pix_638_reg <= Pix_638;
			 Pix_639_reg <= Pix_639;
			 Pix_640_reg <= Pix_640;
			 Pix_641_reg <= Pix_641;
			 Pix_642_reg <= Pix_642;
			 Pix_643_reg <= Pix_643;
			 Pix_644_reg <= Pix_644;
			 Pix_645_reg <= Pix_645;
			 Pix_646_reg <= Pix_646;
			 Pix_647_reg <= Pix_647;
			 Pix_648_reg <= Pix_648;
			 Pix_649_reg <= Pix_649;
			 Pix_650_reg <= Pix_650;
			 Pix_651_reg <= Pix_651;
			 Pix_652_reg <= Pix_652;
			 Pix_653_reg <= Pix_653;
			 Pix_654_reg <= Pix_654;
			 Pix_655_reg <= Pix_655;
			 Pix_656_reg <= Pix_656;
			 Pix_657_reg <= Pix_657;
			 Pix_658_reg <= Pix_658;
			 Pix_659_reg <= Pix_659;
			 Pix_660_reg <= Pix_660;
			 Pix_661_reg <= Pix_661;
			 Pix_662_reg <= Pix_662;
			 Pix_663_reg <= Pix_663;
			 Pix_664_reg <= Pix_664;
			 Pix_665_reg <= Pix_665;
			 Pix_666_reg <= Pix_666;
			 Pix_667_reg <= Pix_667;
			 Pix_668_reg <= Pix_668;
			 Pix_669_reg <= Pix_669;
			 Pix_670_reg <= Pix_670;
			 Pix_671_reg <= Pix_671;
			 Pix_672_reg <= Pix_672;
			 Pix_673_reg <= Pix_673;
			 Pix_674_reg <= Pix_674;
			 Pix_675_reg <= Pix_675;
			 Pix_676_reg <= Pix_676;
			 Pix_677_reg <= Pix_677;
			 Pix_678_reg <= Pix_678;
			 Pix_679_reg <= Pix_679;
			 Pix_680_reg <= Pix_680;
			 Pix_681_reg <= Pix_681;
			 Pix_682_reg <= Pix_682;
			 Pix_683_reg <= Pix_683;
			 Pix_684_reg <= Pix_684;
			 Pix_685_reg <= Pix_685;
			 Pix_686_reg <= Pix_686;
			 Pix_687_reg <= Pix_687;
			 Pix_688_reg <= Pix_688;
			 Pix_689_reg <= Pix_689;
			 Pix_690_reg <= Pix_690;
			 Pix_691_reg <= Pix_691;
			 Pix_692_reg <= Pix_692;
			 Pix_693_reg <= Pix_693;
			 Pix_694_reg <= Pix_694;
			 Pix_695_reg <= Pix_695;
			 Pix_696_reg <= Pix_696;
			 Pix_697_reg <= Pix_697;
			 Pix_698_reg <= Pix_698;
			 Pix_699_reg <= Pix_699;
			 Pix_700_reg <= Pix_700;
			 Pix_701_reg <= Pix_701;
			 Pix_702_reg <= Pix_702;
			 Pix_703_reg <= Pix_703;
			 Pix_704_reg <= Pix_704;
			 Pix_705_reg <= Pix_705;
			 Pix_706_reg <= Pix_706;
			 Pix_707_reg <= Pix_707;
			 Pix_708_reg <= Pix_708;
			 Pix_709_reg <= Pix_709;
			 Pix_710_reg <= Pix_710;
			 Pix_711_reg <= Pix_711;
			 Pix_712_reg <= Pix_712;
			 Pix_713_reg <= Pix_713;
			 Pix_714_reg <= Pix_714;
			 Pix_715_reg <= Pix_715;
			 Pix_716_reg <= Pix_716;
			 Pix_717_reg <= Pix_717;
			 Pix_718_reg <= Pix_718;
			 Pix_719_reg <= Pix_719;
			 Pix_720_reg <= Pix_720;
			 Pix_721_reg <= Pix_721;
			 Pix_722_reg <= Pix_722;
			 Pix_723_reg <= Pix_723;
			 Pix_724_reg <= Pix_724;
			 Pix_725_reg <= Pix_725;
			 Pix_726_reg <= Pix_726;
			 Pix_727_reg <= Pix_727;
			 Pix_728_reg <= Pix_728;
			 Pix_729_reg <= Pix_729;
			 Pix_730_reg <= Pix_730;
			 Pix_731_reg <= Pix_731;
			 Pix_732_reg <= Pix_732;
			 Pix_733_reg <= Pix_733;
			 Pix_734_reg <= Pix_734;
			 Pix_735_reg <= Pix_735;
			 Pix_736_reg <= Pix_736;
			 Pix_737_reg <= Pix_737;
			 Pix_738_reg <= Pix_738;
			 Pix_739_reg <= Pix_739;
			 Pix_740_reg <= Pix_740;
			 Pix_741_reg <= Pix_741;
			 Pix_742_reg <= Pix_742;
			 Pix_743_reg <= Pix_743;
			 Pix_744_reg <= Pix_744;
			 Pix_745_reg <= Pix_745;
			 Pix_746_reg <= Pix_746;
			 Pix_747_reg <= Pix_747;
			 Pix_748_reg <= Pix_748;
			 Pix_749_reg <= Pix_749;
			 Pix_750_reg <= Pix_750;
			 Pix_751_reg <= Pix_751;
			 Pix_752_reg <= Pix_752;
			 Pix_753_reg <= Pix_753;
			 Pix_754_reg <= Pix_754;
			 Pix_755_reg <= Pix_755;
			 Pix_756_reg <= Pix_756;
			 Pix_757_reg <= Pix_757;
			 Pix_758_reg <= Pix_758;
			 Pix_759_reg <= Pix_759;
			 Pix_760_reg <= Pix_760;
			 Pix_761_reg <= Pix_761;
			 Pix_762_reg <= Pix_762;
			 Pix_763_reg <= Pix_763;
			 Pix_764_reg <= Pix_764;
			 Pix_765_reg <= Pix_765;
			 Pix_766_reg <= Pix_766;
			 Pix_767_reg <= Pix_767;
			 Pix_768_reg <= Pix_768;
			 Pix_769_reg <= Pix_769;
			 Pix_770_reg <= Pix_770;
			 Pix_771_reg <= Pix_771;
			 Pix_772_reg <= Pix_772;
			 Pix_773_reg <= Pix_773;
			 Pix_774_reg <= Pix_774;
			 Pix_775_reg <= Pix_775;
			 Pix_776_reg <= Pix_776;
			 Pix_777_reg <= Pix_777;
			 Pix_778_reg <= Pix_778;
			 Pix_779_reg <= Pix_779;
			 Pix_780_reg <= Pix_780;
			 Pix_781_reg <= Pix_781;
			 Pix_782_reg <= Pix_782;
			 Pix_783_reg <= Pix_783;
		end
		else begin
			 Pix_0_reg <= Pix_0_reg;
			 Pix_1_reg <= Pix_1_reg;
			 Pix_2_reg <= Pix_2_reg;
			 Pix_3_reg <= Pix_3_reg;
			 Pix_4_reg <= Pix_4_reg;
			 Pix_5_reg <= Pix_5_reg;
			 Pix_6_reg <= Pix_6_reg;
			 Pix_7_reg <= Pix_7_reg;
			 Pix_8_reg <= Pix_8_reg;
			 Pix_9_reg <= Pix_9_reg;
			 Pix_10_reg <= Pix_10_reg;
			 Pix_11_reg <= Pix_11_reg;
			 Pix_12_reg <= Pix_12_reg;
			 Pix_13_reg <= Pix_13_reg;
			 Pix_14_reg <= Pix_14_reg;
			 Pix_15_reg <= Pix_15_reg;
			 Pix_16_reg <= Pix_16_reg;
			 Pix_17_reg <= Pix_17_reg;
			 Pix_18_reg <= Pix_18_reg;
			 Pix_19_reg <= Pix_19_reg;
			 Pix_20_reg <= Pix_20_reg;
			 Pix_21_reg <= Pix_21_reg;
			 Pix_22_reg <= Pix_22_reg;
			 Pix_23_reg <= Pix_23_reg;
			 Pix_24_reg <= Pix_24_reg;
			 Pix_25_reg <= Pix_25_reg;
			 Pix_26_reg <= Pix_26_reg;
			 Pix_27_reg <= Pix_27_reg;
			 Pix_28_reg <= Pix_28_reg;
			 Pix_29_reg <= Pix_29_reg;
			 Pix_30_reg <= Pix_30_reg;
			 Pix_31_reg <= Pix_31_reg;
			 Pix_32_reg <= Pix_32_reg;
			 Pix_33_reg <= Pix_33_reg;
			 Pix_34_reg <= Pix_34_reg;
			 Pix_35_reg <= Pix_35_reg;
			 Pix_36_reg <= Pix_36_reg;
			 Pix_37_reg <= Pix_37_reg;
			 Pix_38_reg <= Pix_38_reg;
			 Pix_39_reg <= Pix_39_reg;
			 Pix_40_reg <= Pix_40_reg;
			 Pix_41_reg <= Pix_41_reg;
			 Pix_42_reg <= Pix_42_reg;
			 Pix_43_reg <= Pix_43_reg;
			 Pix_44_reg <= Pix_44_reg;
			 Pix_45_reg <= Pix_45_reg;
			 Pix_46_reg <= Pix_46_reg;
			 Pix_47_reg <= Pix_47_reg;
			 Pix_48_reg <= Pix_48_reg;
			 Pix_49_reg <= Pix_49_reg;
			 Pix_50_reg <= Pix_50_reg;
			 Pix_51_reg <= Pix_51_reg;
			 Pix_52_reg <= Pix_52_reg;
			 Pix_53_reg <= Pix_53_reg;
			 Pix_54_reg <= Pix_54_reg;
			 Pix_55_reg <= Pix_55_reg;
			 Pix_56_reg <= Pix_56_reg;
			 Pix_57_reg <= Pix_57_reg;
			 Pix_58_reg <= Pix_58_reg;
			 Pix_59_reg <= Pix_59_reg;
			 Pix_60_reg <= Pix_60_reg;
			 Pix_61_reg <= Pix_61_reg;
			 Pix_62_reg <= Pix_62_reg;
			 Pix_63_reg <= Pix_63_reg;
			 Pix_64_reg <= Pix_64_reg;
			 Pix_65_reg <= Pix_65_reg;
			 Pix_66_reg <= Pix_66_reg;
			 Pix_67_reg <= Pix_67_reg;
			 Pix_68_reg <= Pix_68_reg;
			 Pix_69_reg <= Pix_69_reg;
			 Pix_70_reg <= Pix_70_reg;
			 Pix_71_reg <= Pix_71_reg;
			 Pix_72_reg <= Pix_72_reg;
			 Pix_73_reg <= Pix_73_reg;
			 Pix_74_reg <= Pix_74_reg;
			 Pix_75_reg <= Pix_75_reg;
			 Pix_76_reg <= Pix_76_reg;
			 Pix_77_reg <= Pix_77_reg;
			 Pix_78_reg <= Pix_78_reg;
			 Pix_79_reg <= Pix_79_reg;
			 Pix_80_reg <= Pix_80_reg;
			 Pix_81_reg <= Pix_81_reg;
			 Pix_82_reg <= Pix_82_reg;
			 Pix_83_reg <= Pix_83_reg;
			 Pix_84_reg <= Pix_84_reg;
			 Pix_85_reg <= Pix_85_reg;
			 Pix_86_reg <= Pix_86_reg;
			 Pix_87_reg <= Pix_87_reg;
			 Pix_88_reg <= Pix_88_reg;
			 Pix_89_reg <= Pix_89_reg;
			 Pix_90_reg <= Pix_90_reg;
			 Pix_91_reg <= Pix_91_reg;
			 Pix_92_reg <= Pix_92_reg;
			 Pix_93_reg <= Pix_93_reg;
			 Pix_94_reg <= Pix_94_reg;
			 Pix_95_reg <= Pix_95_reg;
			 Pix_96_reg <= Pix_96_reg;
			 Pix_97_reg <= Pix_97_reg;
			 Pix_98_reg <= Pix_98_reg;
			 Pix_99_reg <= Pix_99_reg;
			 Pix_100_reg <= Pix_100_reg;
			 Pix_101_reg <= Pix_101_reg;
			 Pix_102_reg <= Pix_102_reg;
			 Pix_103_reg <= Pix_103_reg;
			 Pix_104_reg <= Pix_104_reg;
			 Pix_105_reg <= Pix_105_reg;
			 Pix_106_reg <= Pix_106_reg;
			 Pix_107_reg <= Pix_107_reg;
			 Pix_108_reg <= Pix_108_reg;
			 Pix_109_reg <= Pix_109_reg;
			 Pix_110_reg <= Pix_110_reg;
			 Pix_111_reg <= Pix_111_reg;
			 Pix_112_reg <= Pix_112_reg;
			 Pix_113_reg <= Pix_113_reg;
			 Pix_114_reg <= Pix_114_reg;
			 Pix_115_reg <= Pix_115_reg;
			 Pix_116_reg <= Pix_116_reg;
			 Pix_117_reg <= Pix_117_reg;
			 Pix_118_reg <= Pix_118_reg;
			 Pix_119_reg <= Pix_119_reg;
			 Pix_120_reg <= Pix_120_reg;
			 Pix_121_reg <= Pix_121_reg;
			 Pix_122_reg <= Pix_122_reg;
			 Pix_123_reg <= Pix_123_reg;
			 Pix_124_reg <= Pix_124_reg;
			 Pix_125_reg <= Pix_125_reg;
			 Pix_126_reg <= Pix_126_reg;
			 Pix_127_reg <= Pix_127_reg;
			 Pix_128_reg <= Pix_128_reg;
			 Pix_129_reg <= Pix_129_reg;
			 Pix_130_reg <= Pix_130_reg;
			 Pix_131_reg <= Pix_131_reg;
			 Pix_132_reg <= Pix_132_reg;
			 Pix_133_reg <= Pix_133_reg;
			 Pix_134_reg <= Pix_134_reg;
			 Pix_135_reg <= Pix_135_reg;
			 Pix_136_reg <= Pix_136_reg;
			 Pix_137_reg <= Pix_137_reg;
			 Pix_138_reg <= Pix_138_reg;
			 Pix_139_reg <= Pix_139_reg;
			 Pix_140_reg <= Pix_140_reg;
			 Pix_141_reg <= Pix_141_reg;
			 Pix_142_reg <= Pix_142_reg;
			 Pix_143_reg <= Pix_143_reg;
			 Pix_144_reg <= Pix_144_reg;
			 Pix_145_reg <= Pix_145_reg;
			 Pix_146_reg <= Pix_146_reg;
			 Pix_147_reg <= Pix_147_reg;
			 Pix_148_reg <= Pix_148_reg;
			 Pix_149_reg <= Pix_149_reg;
			 Pix_150_reg <= Pix_150_reg;
			 Pix_151_reg <= Pix_151_reg;
			 Pix_152_reg <= Pix_152_reg;
			 Pix_153_reg <= Pix_153_reg;
			 Pix_154_reg <= Pix_154_reg;
			 Pix_155_reg <= Pix_155_reg;
			 Pix_156_reg <= Pix_156_reg;
			 Pix_157_reg <= Pix_157_reg;
			 Pix_158_reg <= Pix_158_reg;
			 Pix_159_reg <= Pix_159_reg;
			 Pix_160_reg <= Pix_160_reg;
			 Pix_161_reg <= Pix_161_reg;
			 Pix_162_reg <= Pix_162_reg;
			 Pix_163_reg <= Pix_163_reg;
			 Pix_164_reg <= Pix_164_reg;
			 Pix_165_reg <= Pix_165_reg;
			 Pix_166_reg <= Pix_166_reg;
			 Pix_167_reg <= Pix_167_reg;
			 Pix_168_reg <= Pix_168_reg;
			 Pix_169_reg <= Pix_169_reg;
			 Pix_170_reg <= Pix_170_reg;
			 Pix_171_reg <= Pix_171_reg;
			 Pix_172_reg <= Pix_172_reg;
			 Pix_173_reg <= Pix_173_reg;
			 Pix_174_reg <= Pix_174_reg;
			 Pix_175_reg <= Pix_175_reg;
			 Pix_176_reg <= Pix_176_reg;
			 Pix_177_reg <= Pix_177_reg;
			 Pix_178_reg <= Pix_178_reg;
			 Pix_179_reg <= Pix_179_reg;
			 Pix_180_reg <= Pix_180_reg;
			 Pix_181_reg <= Pix_181_reg;
			 Pix_182_reg <= Pix_182_reg;
			 Pix_183_reg <= Pix_183_reg;
			 Pix_184_reg <= Pix_184_reg;
			 Pix_185_reg <= Pix_185_reg;
			 Pix_186_reg <= Pix_186_reg;
			 Pix_187_reg <= Pix_187_reg;
			 Pix_188_reg <= Pix_188_reg;
			 Pix_189_reg <= Pix_189_reg;
			 Pix_190_reg <= Pix_190_reg;
			 Pix_191_reg <= Pix_191_reg;
			 Pix_192_reg <= Pix_192_reg;
			 Pix_193_reg <= Pix_193_reg;
			 Pix_194_reg <= Pix_194_reg;
			 Pix_195_reg <= Pix_195_reg;
			 Pix_196_reg <= Pix_196_reg;
			 Pix_197_reg <= Pix_197_reg;
			 Pix_198_reg <= Pix_198_reg;
			 Pix_199_reg <= Pix_199_reg;
			 Pix_200_reg <= Pix_200_reg;
			 Pix_201_reg <= Pix_201_reg;
			 Pix_202_reg <= Pix_202_reg;
			 Pix_203_reg <= Pix_203_reg;
			 Pix_204_reg <= Pix_204_reg;
			 Pix_205_reg <= Pix_205_reg;
			 Pix_206_reg <= Pix_206_reg;
			 Pix_207_reg <= Pix_207_reg;
			 Pix_208_reg <= Pix_208_reg;
			 Pix_209_reg <= Pix_209_reg;
			 Pix_210_reg <= Pix_210_reg;
			 Pix_211_reg <= Pix_211_reg;
			 Pix_212_reg <= Pix_212_reg;
			 Pix_213_reg <= Pix_213_reg;
			 Pix_214_reg <= Pix_214_reg;
			 Pix_215_reg <= Pix_215_reg;
			 Pix_216_reg <= Pix_216_reg;
			 Pix_217_reg <= Pix_217_reg;
			 Pix_218_reg <= Pix_218_reg;
			 Pix_219_reg <= Pix_219_reg;
			 Pix_220_reg <= Pix_220_reg;
			 Pix_221_reg <= Pix_221_reg;
			 Pix_222_reg <= Pix_222_reg;
			 Pix_223_reg <= Pix_223_reg;
			 Pix_224_reg <= Pix_224_reg;
			 Pix_225_reg <= Pix_225_reg;
			 Pix_226_reg <= Pix_226_reg;
			 Pix_227_reg <= Pix_227_reg;
			 Pix_228_reg <= Pix_228_reg;
			 Pix_229_reg <= Pix_229_reg;
			 Pix_230_reg <= Pix_230_reg;
			 Pix_231_reg <= Pix_231_reg;
			 Pix_232_reg <= Pix_232_reg;
			 Pix_233_reg <= Pix_233_reg;
			 Pix_234_reg <= Pix_234_reg;
			 Pix_235_reg <= Pix_235_reg;
			 Pix_236_reg <= Pix_236_reg;
			 Pix_237_reg <= Pix_237_reg;
			 Pix_238_reg <= Pix_238_reg;
			 Pix_239_reg <= Pix_239_reg;
			 Pix_240_reg <= Pix_240_reg;
			 Pix_241_reg <= Pix_241_reg;
			 Pix_242_reg <= Pix_242_reg;
			 Pix_243_reg <= Pix_243_reg;
			 Pix_244_reg <= Pix_244_reg;
			 Pix_245_reg <= Pix_245_reg;
			 Pix_246_reg <= Pix_246_reg;
			 Pix_247_reg <= Pix_247_reg;
			 Pix_248_reg <= Pix_248_reg;
			 Pix_249_reg <= Pix_249_reg;
			 Pix_250_reg <= Pix_250_reg;
			 Pix_251_reg <= Pix_251_reg;
			 Pix_252_reg <= Pix_252_reg;
			 Pix_253_reg <= Pix_253_reg;
			 Pix_254_reg <= Pix_254_reg;
			 Pix_255_reg <= Pix_255_reg;
			 Pix_256_reg <= Pix_256_reg;
			 Pix_257_reg <= Pix_257_reg;
			 Pix_258_reg <= Pix_258_reg;
			 Pix_259_reg <= Pix_259_reg;
			 Pix_260_reg <= Pix_260_reg;
			 Pix_261_reg <= Pix_261_reg;
			 Pix_262_reg <= Pix_262_reg;
			 Pix_263_reg <= Pix_263_reg;
			 Pix_264_reg <= Pix_264_reg;
			 Pix_265_reg <= Pix_265_reg;
			 Pix_266_reg <= Pix_266_reg;
			 Pix_267_reg <= Pix_267_reg;
			 Pix_268_reg <= Pix_268_reg;
			 Pix_269_reg <= Pix_269_reg;
			 Pix_270_reg <= Pix_270_reg;
			 Pix_271_reg <= Pix_271_reg;
			 Pix_272_reg <= Pix_272_reg;
			 Pix_273_reg <= Pix_273_reg;
			 Pix_274_reg <= Pix_274_reg;
			 Pix_275_reg <= Pix_275_reg;
			 Pix_276_reg <= Pix_276_reg;
			 Pix_277_reg <= Pix_277_reg;
			 Pix_278_reg <= Pix_278_reg;
			 Pix_279_reg <= Pix_279_reg;
			 Pix_280_reg <= Pix_280_reg;
			 Pix_281_reg <= Pix_281_reg;
			 Pix_282_reg <= Pix_282_reg;
			 Pix_283_reg <= Pix_283_reg;
			 Pix_284_reg <= Pix_284_reg;
			 Pix_285_reg <= Pix_285_reg;
			 Pix_286_reg <= Pix_286_reg;
			 Pix_287_reg <= Pix_287_reg;
			 Pix_288_reg <= Pix_288_reg;
			 Pix_289_reg <= Pix_289_reg;
			 Pix_290_reg <= Pix_290_reg;
			 Pix_291_reg <= Pix_291_reg;
			 Pix_292_reg <= Pix_292_reg;
			 Pix_293_reg <= Pix_293_reg;
			 Pix_294_reg <= Pix_294_reg;
			 Pix_295_reg <= Pix_295_reg;
			 Pix_296_reg <= Pix_296_reg;
			 Pix_297_reg <= Pix_297_reg;
			 Pix_298_reg <= Pix_298_reg;
			 Pix_299_reg <= Pix_299_reg;
			 Pix_300_reg <= Pix_300_reg;
			 Pix_301_reg <= Pix_301_reg;
			 Pix_302_reg <= Pix_302_reg;
			 Pix_303_reg <= Pix_303_reg;
			 Pix_304_reg <= Pix_304_reg;
			 Pix_305_reg <= Pix_305_reg;
			 Pix_306_reg <= Pix_306_reg;
			 Pix_307_reg <= Pix_307_reg;
			 Pix_308_reg <= Pix_308_reg;
			 Pix_309_reg <= Pix_309_reg;
			 Pix_310_reg <= Pix_310_reg;
			 Pix_311_reg <= Pix_311_reg;
			 Pix_312_reg <= Pix_312_reg;
			 Pix_313_reg <= Pix_313_reg;
			 Pix_314_reg <= Pix_314_reg;
			 Pix_315_reg <= Pix_315_reg;
			 Pix_316_reg <= Pix_316_reg;
			 Pix_317_reg <= Pix_317_reg;
			 Pix_318_reg <= Pix_318_reg;
			 Pix_319_reg <= Pix_319_reg;
			 Pix_320_reg <= Pix_320_reg;
			 Pix_321_reg <= Pix_321_reg;
			 Pix_322_reg <= Pix_322_reg;
			 Pix_323_reg <= Pix_323_reg;
			 Pix_324_reg <= Pix_324_reg;
			 Pix_325_reg <= Pix_325_reg;
			 Pix_326_reg <= Pix_326_reg;
			 Pix_327_reg <= Pix_327_reg;
			 Pix_328_reg <= Pix_328_reg;
			 Pix_329_reg <= Pix_329_reg;
			 Pix_330_reg <= Pix_330_reg;
			 Pix_331_reg <= Pix_331_reg;
			 Pix_332_reg <= Pix_332_reg;
			 Pix_333_reg <= Pix_333_reg;
			 Pix_334_reg <= Pix_334_reg;
			 Pix_335_reg <= Pix_335_reg;
			 Pix_336_reg <= Pix_336_reg;
			 Pix_337_reg <= Pix_337_reg;
			 Pix_338_reg <= Pix_338_reg;
			 Pix_339_reg <= Pix_339_reg;
			 Pix_340_reg <= Pix_340_reg;
			 Pix_341_reg <= Pix_341_reg;
			 Pix_342_reg <= Pix_342_reg;
			 Pix_343_reg <= Pix_343_reg;
			 Pix_344_reg <= Pix_344_reg;
			 Pix_345_reg <= Pix_345_reg;
			 Pix_346_reg <= Pix_346_reg;
			 Pix_347_reg <= Pix_347_reg;
			 Pix_348_reg <= Pix_348_reg;
			 Pix_349_reg <= Pix_349_reg;
			 Pix_350_reg <= Pix_350_reg;
			 Pix_351_reg <= Pix_351_reg;
			 Pix_352_reg <= Pix_352_reg;
			 Pix_353_reg <= Pix_353_reg;
			 Pix_354_reg <= Pix_354_reg;
			 Pix_355_reg <= Pix_355_reg;
			 Pix_356_reg <= Pix_356_reg;
			 Pix_357_reg <= Pix_357_reg;
			 Pix_358_reg <= Pix_358_reg;
			 Pix_359_reg <= Pix_359_reg;
			 Pix_360_reg <= Pix_360_reg;
			 Pix_361_reg <= Pix_361_reg;
			 Pix_362_reg <= Pix_362_reg;
			 Pix_363_reg <= Pix_363_reg;
			 Pix_364_reg <= Pix_364_reg;
			 Pix_365_reg <= Pix_365_reg;
			 Pix_366_reg <= Pix_366_reg;
			 Pix_367_reg <= Pix_367_reg;
			 Pix_368_reg <= Pix_368_reg;
			 Pix_369_reg <= Pix_369_reg;
			 Pix_370_reg <= Pix_370_reg;
			 Pix_371_reg <= Pix_371_reg;
			 Pix_372_reg <= Pix_372_reg;
			 Pix_373_reg <= Pix_373_reg;
			 Pix_374_reg <= Pix_374_reg;
			 Pix_375_reg <= Pix_375_reg;
			 Pix_376_reg <= Pix_376_reg;
			 Pix_377_reg <= Pix_377_reg;
			 Pix_378_reg <= Pix_378_reg;
			 Pix_379_reg <= Pix_379_reg;
			 Pix_380_reg <= Pix_380_reg;
			 Pix_381_reg <= Pix_381_reg;
			 Pix_382_reg <= Pix_382_reg;
			 Pix_383_reg <= Pix_383_reg;
			 Pix_384_reg <= Pix_384_reg;
			 Pix_385_reg <= Pix_385_reg;
			 Pix_386_reg <= Pix_386_reg;
			 Pix_387_reg <= Pix_387_reg;
			 Pix_388_reg <= Pix_388_reg;
			 Pix_389_reg <= Pix_389_reg;
			 Pix_390_reg <= Pix_390_reg;
			 Pix_391_reg <= Pix_391_reg;
			 Pix_392_reg <= Pix_392_reg;
			 Pix_393_reg <= Pix_393_reg;
			 Pix_394_reg <= Pix_394_reg;
			 Pix_395_reg <= Pix_395_reg;
			 Pix_396_reg <= Pix_396_reg;
			 Pix_397_reg <= Pix_397_reg;
			 Pix_398_reg <= Pix_398_reg;
			 Pix_399_reg <= Pix_399_reg;
			 Pix_400_reg <= Pix_400_reg;
			 Pix_401_reg <= Pix_401_reg;
			 Pix_402_reg <= Pix_402_reg;
			 Pix_403_reg <= Pix_403_reg;
			 Pix_404_reg <= Pix_404_reg;
			 Pix_405_reg <= Pix_405_reg;
			 Pix_406_reg <= Pix_406_reg;
			 Pix_407_reg <= Pix_407_reg;
			 Pix_408_reg <= Pix_408_reg;
			 Pix_409_reg <= Pix_409_reg;
			 Pix_410_reg <= Pix_410_reg;
			 Pix_411_reg <= Pix_411_reg;
			 Pix_412_reg <= Pix_412_reg;
			 Pix_413_reg <= Pix_413_reg;
			 Pix_414_reg <= Pix_414_reg;
			 Pix_415_reg <= Pix_415_reg;
			 Pix_416_reg <= Pix_416_reg;
			 Pix_417_reg <= Pix_417_reg;
			 Pix_418_reg <= Pix_418_reg;
			 Pix_419_reg <= Pix_419_reg;
			 Pix_420_reg <= Pix_420_reg;
			 Pix_421_reg <= Pix_421_reg;
			 Pix_422_reg <= Pix_422_reg;
			 Pix_423_reg <= Pix_423_reg;
			 Pix_424_reg <= Pix_424_reg;
			 Pix_425_reg <= Pix_425_reg;
			 Pix_426_reg <= Pix_426_reg;
			 Pix_427_reg <= Pix_427_reg;
			 Pix_428_reg <= Pix_428_reg;
			 Pix_429_reg <= Pix_429_reg;
			 Pix_430_reg <= Pix_430_reg;
			 Pix_431_reg <= Pix_431_reg;
			 Pix_432_reg <= Pix_432_reg;
			 Pix_433_reg <= Pix_433_reg;
			 Pix_434_reg <= Pix_434_reg;
			 Pix_435_reg <= Pix_435_reg;
			 Pix_436_reg <= Pix_436_reg;
			 Pix_437_reg <= Pix_437_reg;
			 Pix_438_reg <= Pix_438_reg;
			 Pix_439_reg <= Pix_439_reg;
			 Pix_440_reg <= Pix_440_reg;
			 Pix_441_reg <= Pix_441_reg;
			 Pix_442_reg <= Pix_442_reg;
			 Pix_443_reg <= Pix_443_reg;
			 Pix_444_reg <= Pix_444_reg;
			 Pix_445_reg <= Pix_445_reg;
			 Pix_446_reg <= Pix_446_reg;
			 Pix_447_reg <= Pix_447_reg;
			 Pix_448_reg <= Pix_448_reg;
			 Pix_449_reg <= Pix_449_reg;
			 Pix_450_reg <= Pix_450_reg;
			 Pix_451_reg <= Pix_451_reg;
			 Pix_452_reg <= Pix_452_reg;
			 Pix_453_reg <= Pix_453_reg;
			 Pix_454_reg <= Pix_454_reg;
			 Pix_455_reg <= Pix_455_reg;
			 Pix_456_reg <= Pix_456_reg;
			 Pix_457_reg <= Pix_457_reg;
			 Pix_458_reg <= Pix_458_reg;
			 Pix_459_reg <= Pix_459_reg;
			 Pix_460_reg <= Pix_460_reg;
			 Pix_461_reg <= Pix_461_reg;
			 Pix_462_reg <= Pix_462_reg;
			 Pix_463_reg <= Pix_463_reg;
			 Pix_464_reg <= Pix_464_reg;
			 Pix_465_reg <= Pix_465_reg;
			 Pix_466_reg <= Pix_466_reg;
			 Pix_467_reg <= Pix_467_reg;
			 Pix_468_reg <= Pix_468_reg;
			 Pix_469_reg <= Pix_469_reg;
			 Pix_470_reg <= Pix_470_reg;
			 Pix_471_reg <= Pix_471_reg;
			 Pix_472_reg <= Pix_472_reg;
			 Pix_473_reg <= Pix_473_reg;
			 Pix_474_reg <= Pix_474_reg;
			 Pix_475_reg <= Pix_475_reg;
			 Pix_476_reg <= Pix_476_reg;
			 Pix_477_reg <= Pix_477_reg;
			 Pix_478_reg <= Pix_478_reg;
			 Pix_479_reg <= Pix_479_reg;
			 Pix_480_reg <= Pix_480_reg;
			 Pix_481_reg <= Pix_481_reg;
			 Pix_482_reg <= Pix_482_reg;
			 Pix_483_reg <= Pix_483_reg;
			 Pix_484_reg <= Pix_484_reg;
			 Pix_485_reg <= Pix_485_reg;
			 Pix_486_reg <= Pix_486_reg;
			 Pix_487_reg <= Pix_487_reg;
			 Pix_488_reg <= Pix_488_reg;
			 Pix_489_reg <= Pix_489_reg;
			 Pix_490_reg <= Pix_490_reg;
			 Pix_491_reg <= Pix_491_reg;
			 Pix_492_reg <= Pix_492_reg;
			 Pix_493_reg <= Pix_493_reg;
			 Pix_494_reg <= Pix_494_reg;
			 Pix_495_reg <= Pix_495_reg;
			 Pix_496_reg <= Pix_496_reg;
			 Pix_497_reg <= Pix_497_reg;
			 Pix_498_reg <= Pix_498_reg;
			 Pix_499_reg <= Pix_499_reg;
			 Pix_500_reg <= Pix_500_reg;
			 Pix_501_reg <= Pix_501_reg;
			 Pix_502_reg <= Pix_502_reg;
			 Pix_503_reg <= Pix_503_reg;
			 Pix_504_reg <= Pix_504_reg;
			 Pix_505_reg <= Pix_505_reg;
			 Pix_506_reg <= Pix_506_reg;
			 Pix_507_reg <= Pix_507_reg;
			 Pix_508_reg <= Pix_508_reg;
			 Pix_509_reg <= Pix_509_reg;
			 Pix_510_reg <= Pix_510_reg;
			 Pix_511_reg <= Pix_511_reg;
			 Pix_512_reg <= Pix_512_reg;
			 Pix_513_reg <= Pix_513_reg;
			 Pix_514_reg <= Pix_514_reg;
			 Pix_515_reg <= Pix_515_reg;
			 Pix_516_reg <= Pix_516_reg;
			 Pix_517_reg <= Pix_517_reg;
			 Pix_518_reg <= Pix_518_reg;
			 Pix_519_reg <= Pix_519_reg;
			 Pix_520_reg <= Pix_520_reg;
			 Pix_521_reg <= Pix_521_reg;
			 Pix_522_reg <= Pix_522_reg;
			 Pix_523_reg <= Pix_523_reg;
			 Pix_524_reg <= Pix_524_reg;
			 Pix_525_reg <= Pix_525_reg;
			 Pix_526_reg <= Pix_526_reg;
			 Pix_527_reg <= Pix_527_reg;
			 Pix_528_reg <= Pix_528_reg;
			 Pix_529_reg <= Pix_529_reg;
			 Pix_530_reg <= Pix_530_reg;
			 Pix_531_reg <= Pix_531_reg;
			 Pix_532_reg <= Pix_532_reg;
			 Pix_533_reg <= Pix_533_reg;
			 Pix_534_reg <= Pix_534_reg;
			 Pix_535_reg <= Pix_535_reg;
			 Pix_536_reg <= Pix_536_reg;
			 Pix_537_reg <= Pix_537_reg;
			 Pix_538_reg <= Pix_538_reg;
			 Pix_539_reg <= Pix_539_reg;
			 Pix_540_reg <= Pix_540_reg;
			 Pix_541_reg <= Pix_541_reg;
			 Pix_542_reg <= Pix_542_reg;
			 Pix_543_reg <= Pix_543_reg;
			 Pix_544_reg <= Pix_544_reg;
			 Pix_545_reg <= Pix_545_reg;
			 Pix_546_reg <= Pix_546_reg;
			 Pix_547_reg <= Pix_547_reg;
			 Pix_548_reg <= Pix_548_reg;
			 Pix_549_reg <= Pix_549_reg;
			 Pix_550_reg <= Pix_550_reg;
			 Pix_551_reg <= Pix_551_reg;
			 Pix_552_reg <= Pix_552_reg;
			 Pix_553_reg <= Pix_553_reg;
			 Pix_554_reg <= Pix_554_reg;
			 Pix_555_reg <= Pix_555_reg;
			 Pix_556_reg <= Pix_556_reg;
			 Pix_557_reg <= Pix_557_reg;
			 Pix_558_reg <= Pix_558_reg;
			 Pix_559_reg <= Pix_559_reg;
			 Pix_560_reg <= Pix_560_reg;
			 Pix_561_reg <= Pix_561_reg;
			 Pix_562_reg <= Pix_562_reg;
			 Pix_563_reg <= Pix_563_reg;
			 Pix_564_reg <= Pix_564_reg;
			 Pix_565_reg <= Pix_565_reg;
			 Pix_566_reg <= Pix_566_reg;
			 Pix_567_reg <= Pix_567_reg;
			 Pix_568_reg <= Pix_568_reg;
			 Pix_569_reg <= Pix_569_reg;
			 Pix_570_reg <= Pix_570_reg;
			 Pix_571_reg <= Pix_571_reg;
			 Pix_572_reg <= Pix_572_reg;
			 Pix_573_reg <= Pix_573_reg;
			 Pix_574_reg <= Pix_574_reg;
			 Pix_575_reg <= Pix_575_reg;
			 Pix_576_reg <= Pix_576_reg;
			 Pix_577_reg <= Pix_577_reg;
			 Pix_578_reg <= Pix_578_reg;
			 Pix_579_reg <= Pix_579_reg;
			 Pix_580_reg <= Pix_580_reg;
			 Pix_581_reg <= Pix_581_reg;
			 Pix_582_reg <= Pix_582_reg;
			 Pix_583_reg <= Pix_583_reg;
			 Pix_584_reg <= Pix_584_reg;
			 Pix_585_reg <= Pix_585_reg;
			 Pix_586_reg <= Pix_586_reg;
			 Pix_587_reg <= Pix_587_reg;
			 Pix_588_reg <= Pix_588_reg;
			 Pix_589_reg <= Pix_589_reg;
			 Pix_590_reg <= Pix_590_reg;
			 Pix_591_reg <= Pix_591_reg;
			 Pix_592_reg <= Pix_592_reg;
			 Pix_593_reg <= Pix_593_reg;
			 Pix_594_reg <= Pix_594_reg;
			 Pix_595_reg <= Pix_595_reg;
			 Pix_596_reg <= Pix_596_reg;
			 Pix_597_reg <= Pix_597_reg;
			 Pix_598_reg <= Pix_598_reg;
			 Pix_599_reg <= Pix_599_reg;
			 Pix_600_reg <= Pix_600_reg;
			 Pix_601_reg <= Pix_601_reg;
			 Pix_602_reg <= Pix_602_reg;
			 Pix_603_reg <= Pix_603_reg;
			 Pix_604_reg <= Pix_604_reg;
			 Pix_605_reg <= Pix_605_reg;
			 Pix_606_reg <= Pix_606_reg;
			 Pix_607_reg <= Pix_607_reg;
			 Pix_608_reg <= Pix_608_reg;
			 Pix_609_reg <= Pix_609_reg;
			 Pix_610_reg <= Pix_610_reg;
			 Pix_611_reg <= Pix_611_reg;
			 Pix_612_reg <= Pix_612_reg;
			 Pix_613_reg <= Pix_613_reg;
			 Pix_614_reg <= Pix_614_reg;
			 Pix_615_reg <= Pix_615_reg;
			 Pix_616_reg <= Pix_616_reg;
			 Pix_617_reg <= Pix_617_reg;
			 Pix_618_reg <= Pix_618_reg;
			 Pix_619_reg <= Pix_619_reg;
			 Pix_620_reg <= Pix_620_reg;
			 Pix_621_reg <= Pix_621_reg;
			 Pix_622_reg <= Pix_622_reg;
			 Pix_623_reg <= Pix_623_reg;
			 Pix_624_reg <= Pix_624_reg;
			 Pix_625_reg <= Pix_625_reg;
			 Pix_626_reg <= Pix_626_reg;
			 Pix_627_reg <= Pix_627_reg;
			 Pix_628_reg <= Pix_628_reg;
			 Pix_629_reg <= Pix_629_reg;
			 Pix_630_reg <= Pix_630_reg;
			 Pix_631_reg <= Pix_631_reg;
			 Pix_632_reg <= Pix_632_reg;
			 Pix_633_reg <= Pix_633_reg;
			 Pix_634_reg <= Pix_634_reg;
			 Pix_635_reg <= Pix_635_reg;
			 Pix_636_reg <= Pix_636_reg;
			 Pix_637_reg <= Pix_637_reg;
			 Pix_638_reg <= Pix_638_reg;
			 Pix_639_reg <= Pix_639_reg;
			 Pix_640_reg <= Pix_640_reg;
			 Pix_641_reg <= Pix_641_reg;
			 Pix_642_reg <= Pix_642_reg;
			 Pix_643_reg <= Pix_643_reg;
			 Pix_644_reg <= Pix_644_reg;
			 Pix_645_reg <= Pix_645_reg;
			 Pix_646_reg <= Pix_646_reg;
			 Pix_647_reg <= Pix_647_reg;
			 Pix_648_reg <= Pix_648_reg;
			 Pix_649_reg <= Pix_649_reg;
			 Pix_650_reg <= Pix_650_reg;
			 Pix_651_reg <= Pix_651_reg;
			 Pix_652_reg <= Pix_652_reg;
			 Pix_653_reg <= Pix_653_reg;
			 Pix_654_reg <= Pix_654_reg;
			 Pix_655_reg <= Pix_655_reg;
			 Pix_656_reg <= Pix_656_reg;
			 Pix_657_reg <= Pix_657_reg;
			 Pix_658_reg <= Pix_658_reg;
			 Pix_659_reg <= Pix_659_reg;
			 Pix_660_reg <= Pix_660_reg;
			 Pix_661_reg <= Pix_661_reg;
			 Pix_662_reg <= Pix_662_reg;
			 Pix_663_reg <= Pix_663_reg;
			 Pix_664_reg <= Pix_664_reg;
			 Pix_665_reg <= Pix_665_reg;
			 Pix_666_reg <= Pix_666_reg;
			 Pix_667_reg <= Pix_667_reg;
			 Pix_668_reg <= Pix_668_reg;
			 Pix_669_reg <= Pix_669_reg;
			 Pix_670_reg <= Pix_670_reg;
			 Pix_671_reg <= Pix_671_reg;
			 Pix_672_reg <= Pix_672_reg;
			 Pix_673_reg <= Pix_673_reg;
			 Pix_674_reg <= Pix_674_reg;
			 Pix_675_reg <= Pix_675_reg;
			 Pix_676_reg <= Pix_676_reg;
			 Pix_677_reg <= Pix_677_reg;
			 Pix_678_reg <= Pix_678_reg;
			 Pix_679_reg <= Pix_679_reg;
			 Pix_680_reg <= Pix_680_reg;
			 Pix_681_reg <= Pix_681_reg;
			 Pix_682_reg <= Pix_682_reg;
			 Pix_683_reg <= Pix_683_reg;
			 Pix_684_reg <= Pix_684_reg;
			 Pix_685_reg <= Pix_685_reg;
			 Pix_686_reg <= Pix_686_reg;
			 Pix_687_reg <= Pix_687_reg;
			 Pix_688_reg <= Pix_688_reg;
			 Pix_689_reg <= Pix_689_reg;
			 Pix_690_reg <= Pix_690_reg;
			 Pix_691_reg <= Pix_691_reg;
			 Pix_692_reg <= Pix_692_reg;
			 Pix_693_reg <= Pix_693_reg;
			 Pix_694_reg <= Pix_694_reg;
			 Pix_695_reg <= Pix_695_reg;
			 Pix_696_reg <= Pix_696_reg;
			 Pix_697_reg <= Pix_697_reg;
			 Pix_698_reg <= Pix_698_reg;
			 Pix_699_reg <= Pix_699_reg;
			 Pix_700_reg <= Pix_700_reg;
			 Pix_701_reg <= Pix_701_reg;
			 Pix_702_reg <= Pix_702_reg;
			 Pix_703_reg <= Pix_703_reg;
			 Pix_704_reg <= Pix_704_reg;
			 Pix_705_reg <= Pix_705_reg;
			 Pix_706_reg <= Pix_706_reg;
			 Pix_707_reg <= Pix_707_reg;
			 Pix_708_reg <= Pix_708_reg;
			 Pix_709_reg <= Pix_709_reg;
			 Pix_710_reg <= Pix_710_reg;
			 Pix_711_reg <= Pix_711_reg;
			 Pix_712_reg <= Pix_712_reg;
			 Pix_713_reg <= Pix_713_reg;
			 Pix_714_reg <= Pix_714_reg;
			 Pix_715_reg <= Pix_715_reg;
			 Pix_716_reg <= Pix_716_reg;
			 Pix_717_reg <= Pix_717_reg;
			 Pix_718_reg <= Pix_718_reg;
			 Pix_719_reg <= Pix_719_reg;
			 Pix_720_reg <= Pix_720_reg;
			 Pix_721_reg <= Pix_721_reg;
			 Pix_722_reg <= Pix_722_reg;
			 Pix_723_reg <= Pix_723_reg;
			 Pix_724_reg <= Pix_724_reg;
			 Pix_725_reg <= Pix_725_reg;
			 Pix_726_reg <= Pix_726_reg;
			 Pix_727_reg <= Pix_727_reg;
			 Pix_728_reg <= Pix_728_reg;
			 Pix_729_reg <= Pix_729_reg;
			 Pix_730_reg <= Pix_730_reg;
			 Pix_731_reg <= Pix_731_reg;
			 Pix_732_reg <= Pix_732_reg;
			 Pix_733_reg <= Pix_733_reg;
			 Pix_734_reg <= Pix_734_reg;
			 Pix_735_reg <= Pix_735_reg;
			 Pix_736_reg <= Pix_736_reg;
			 Pix_737_reg <= Pix_737_reg;
			 Pix_738_reg <= Pix_738_reg;
			 Pix_739_reg <= Pix_739_reg;
			 Pix_740_reg <= Pix_740_reg;
			 Pix_741_reg <= Pix_741_reg;
			 Pix_742_reg <= Pix_742_reg;
			 Pix_743_reg <= Pix_743_reg;
			 Pix_744_reg <= Pix_744_reg;
			 Pix_745_reg <= Pix_745_reg;
			 Pix_746_reg <= Pix_746_reg;
			 Pix_747_reg <= Pix_747_reg;
			 Pix_748_reg <= Pix_748_reg;
			 Pix_749_reg <= Pix_749_reg;
			 Pix_750_reg <= Pix_750_reg;
			 Pix_751_reg <= Pix_751_reg;
			 Pix_752_reg <= Pix_752_reg;
			 Pix_753_reg <= Pix_753_reg;
			 Pix_754_reg <= Pix_754_reg;
			 Pix_755_reg <= Pix_755_reg;
			 Pix_756_reg <= Pix_756_reg;
			 Pix_757_reg <= Pix_757_reg;
			 Pix_758_reg <= Pix_758_reg;
			 Pix_759_reg <= Pix_759_reg;
			 Pix_760_reg <= Pix_760_reg;
			 Pix_761_reg <= Pix_761_reg;
			 Pix_762_reg <= Pix_762_reg;
			 Pix_763_reg <= Pix_763_reg;
			 Pix_764_reg <= Pix_764_reg;
			 Pix_765_reg <= Pix_765_reg;
			 Pix_766_reg <= Pix_766_reg;
			 Pix_767_reg <= Pix_767_reg;
			 Pix_768_reg <= Pix_768_reg;
			 Pix_769_reg <= Pix_769_reg;
			 Pix_770_reg <= Pix_770_reg;
			 Pix_771_reg <= Pix_771_reg;
			 Pix_772_reg <= Pix_772_reg;
			 Pix_773_reg <= Pix_773_reg;
			 Pix_774_reg <= Pix_774_reg;
			 Pix_775_reg <= Pix_775_reg;
			 Pix_776_reg <= Pix_776_reg;
			 Pix_777_reg <= Pix_777_reg;
			 Pix_778_reg <= Pix_778_reg;
			 Pix_779_reg <= Pix_779_reg;
			 Pix_780_reg <= Pix_780_reg;
			 Pix_781_reg <= Pix_781_reg;
			 Pix_782_reg <= Pix_782_reg;
			 Pix_783_reg <= Pix_783_reg;
		end
	end
endmodule
	